CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
5 4 0.500000 0.500000
176 79 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
28
5 4081~
219 800 78 0 3 22
0 10 4 3
0
0 0 624 180
4 4081
-7 -24 21 -16
4 U11A
-16 -25 12 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
5130 0 0
2
42185.9 0
0
9 Inverter~
13 847 158 0 2 22
0 16 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
391 0 0
2
42185.9 0
0
5 4012~
219 982 98 0 5 22
0 15 14 13 12 11
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 4 0
1 U
3124 0 0
2
42185.9 0
0
5 4071~
219 887 45 0 3 22
0 11 2 4
0
0 0 624 180
4 4071
-7 -24 21 -16
3 U9A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3421 0 0
2
42185.9 0
0
9 Inverter~
13 1051 237 0 2 22
0 6 5
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
8157 0 0
2
42185.9 0
0
5 4011~
219 1107 228 0 3 22
0 7 5 2
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
42185.9 0
0
9 Inverter~
13 831 238 0 2 22
0 13 18
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
8901 0 0
2
42185.9 0
0
9 Inverter~
13 830 215 0 2 22
0 17 14
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
7361 0 0
2
42185.8 0
0
5 4012~
219 885 219 0 5 22
0 16 14 18 12 10
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 4 0
1 U
4747 0 0
2
42185.8 0
0
9 Inverter~
13 588 191 0 2 22
0 26 27
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U12C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
972 0 0
2
42185.8 0
0
9 Inverter~
13 589 231 0 2 22
0 24 29
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3472 0 0
2
42185.8 0
0
5 4012~
219 643 226 0 5 22
0 27 25 29 23 28
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 1 0
1 U
9998 0 0
2
42185.8 0
0
2 +V
167 928 118 0 1 3
0 30
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3536 0 0
2
42185.8 0
0
2 +V
167 707 123 0 1 3
0 31
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4597 0 0
2
42185.8 0
0
2 +V
167 460 126 0 1 3
0 32
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3835 0 0
2
42185.8 0
0
9 Inverter~
13 340 251 0 2 22
0 20 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3670 0 0
2
42185.8 0
0
9 Inverter~
13 342 225 0 2 22
0 21 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
5616 0 0
2
42185.8 0
0
5 4012~
219 391 229 0 5 22
0 22 35 34 19 33
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 1 0
1 U
9323 0 0
2
42185.8 0
0
12 Hex Display~
7 153 439 0 16 19
10 6 7 8 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
317 0 0
2
42185.8 0
0
12 Hex Display~
7 188 439 0 16 19
10 12 13 17 16 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3108 0 0
2
42185.8 0
0
12 Hex Display~
7 231 439 0 18 19
10 23 24 25 26 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4299 0 0
2
42185.8 0
0
12 Hex Display~
7 266 439 0 18 19
10 19 20 21 22 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9672 0 0
2
42185.8 0
0
2 +V
167 169 121 0 1 3
0 36
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7876 0 0
2
42185.8 0
0
7 Pulser~
4 74 207 0 10 12
0 38 39 37 40 0 0 5 5 5
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6369 0 0
2
42185.8 0
0
7 74LS163
126 985 198 0 14 29
0 30 30 3 30 41 42 43 44 2
45 9 8 7 6
0
0 0 4848 0
8 74LS163A
-28 -51 28 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
9172 0 0
2
42185.8 0
0
7 74LS163
126 764 199 0 14 29
0 31 31 28 31 46 47 48 49 3
50 16 17 13 12
0
0 0 4848 0
8 74LS163A
-28 -51 28 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
7100 0 0
2
42185.8 0
0
7 74LS163
126 508 204 0 14 29
0 32 32 33 32 51 52 53 54 28
55 26 25 24 23
0
0 0 4848 0
8 74LS163A
-28 -51 28 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
3820 0 0
2
42185.8 0
0
7 74LS163
126 246 207 0 14 29
0 36 36 37 36 56 57 58 59 33
60 22 21 20 19
0
0 0 4848 0
8 74LS163A
-28 -51 28 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
7678 0 0
2
42185.8 0
0
67
9 0 2 0 0 4096 0 25 0 0 14 2
1023 171
1134 171
3 0 3 0 0 12416 0 25 0 0 3 4
953 189
876 189
876 104
752 104
3 9 3 0 0 0 0 1 26 0 0 5
773 78
752 78
752 127
802 127
802 172
3 2 4 0 0 4224 0 4 1 0 0 4
860 45
822 45
822 69
818 69
2 2 5 0 0 4224 0 5 6 0 0 2
1072 237
1083 237
0 1 6 0 0 8192 0 0 5 7 0 3
1027 239
1027 237
1036 237
14 0 6 0 0 8192 0 25 0 0 8 3
1017 234
1027 234
1027 271
0 1 6 0 0 8320 0 0 19 0 0 4
1027 268
1027 576
162 576
162 463
0 2 7 0 0 8320 0 0 19 20 0 4
1032 225
1032 589
156 589
156 463
12 3 8 0 0 12416 0 25 19 0 0 5
1017 216
1067 216
1067 598
150 598
150 463
11 4 9 0 0 12416 0 25 19 0 0 5
1017 207
1157 207
1157 610
144 610
144 463
5 1 10 0 0 8320 0 9 1 0 0 6
912 219
918 219
918 127
856 127
856 87
818 87
1 5 11 0 0 4224 0 4 3 0 0 4
906 54
1057 54
1057 98
1009 98
3 2 2 0 0 8320 0 6 4 0 0 3
1134 228
1134 36
906 36
0 4 12 0 0 8192 0 0 3 26 0 4
859 260
946 260
946 112
958 112
0 3 13 0 0 12288 0 0 3 23 0 5
776 523
776 395
940 395
940 103
958 103
0 2 14 0 0 12416 0 0 3 29 0 5
854 215
854 175
899 175
899 94
958 94
2 1 15 0 0 8320 0 2 3 0 0 4
868 158
887 158
887 85
958 85
0 1 16 0 0 4096 0 0 2 21 0 5
814 206
814 181
826 181
826 158
832 158
13 1 7 0 0 0 0 25 6 0 0 4
1017 225
1075 225
1075 219
1083 219
0 4 16 0 0 8320 0 0 20 25 0 4
814 206
814 556
179 556
179 463
0 3 17 0 0 8320 0 0 20 30 0 4
806 217
806 533
185 533
185 463
0 2 13 0 0 8320 0 0 20 28 0 4
803 226
803 523
191 523
191 463
0 1 12 0 0 8320 0 0 20 26 0 4
796 260
796 510
197 510
197 463
11 1 16 0 0 0 0 26 9 0 0 3
796 208
796 206
861 206
14 4 12 0 0 0 0 26 9 0 0 4
796 235
796 260
861 260
861 233
2 3 18 0 0 4224 0 7 9 0 0 3
852 238
852 224
861 224
1 13 13 0 0 0 0 7 26 0 0 4
816 238
810 238
810 226
796 226
2 2 14 0 0 0 0 8 9 0 0 2
851 215
861 215
12 1 17 0 0 0 0 26 8 0 0 4
796 217
807 217
807 215
815 215
0 1 19 0 0 4224 0 0 22 58 0 3
286 243
286 463
275 463
0 2 20 0 0 4224 0 0 22 60 0 4
290 234
290 488
269 488
269 463
0 3 21 0 0 4224 0 0 22 62 0 4
302 225
302 483
263 483
263 463
0 4 22 0 0 4224 0 0 22 63 0 4
312 216
312 478
257 478
257 463
0 1 23 0 0 8320 0 0 21 43 0 4
569 240
569 496
240 496
240 463
0 2 24 0 0 24704 0 0 21 45 0 8
547 231
547 153
614 153
614 422
622 422
622 486
234 486
234 463
0 3 25 0 0 8320 0 0 21 44 0 4
552 222
552 491
228 491
228 463
0 4 26 0 0 16512 0 0 21 40 0 6
548 213
548 158
558 158
558 486
222 486
222 463
2 1 27 0 0 8320 0 10 12 0 0 4
609 191
613 191
613 213
619 213
11 1 26 0 0 0 0 27 10 0 0 4
540 213
565 213
565 191
573 191
3 0 28 0 0 4096 0 26 0 0 42 2
732 190
689 190
9 5 28 0 0 4224 0 27 12 0 0 4
546 177
689 177
689 226
670 226
14 4 23 0 0 0 0 27 12 0 0 6
540 240
570 240
570 243
614 243
614 240
619 240
12 2 25 0 0 0 0 27 12 0 0 6
540 222
574 222
574 208
605 208
605 222
619 222
13 1 24 0 0 0 0 27 11 0 0 2
540 231
574 231
2 3 29 0 0 4224 0 11 12 0 0 2
610 231
619 231
1 0 30 0 0 4096 0 25 0 0 49 2
953 171
928 171
2 0 30 0 0 0 0 25 0 0 49 2
953 180
928 180
1 4 30 0 0 4224 0 13 25 0 0 3
928 127
928 198
947 198
1 0 31 0 0 4096 0 26 0 0 52 2
732 172
707 172
2 0 31 0 0 0 0 26 0 0 52 2
732 181
707 181
1 4 31 0 0 4224 0 14 26 0 0 3
707 132
707 199
726 199
1 0 32 0 0 4096 0 27 0 0 55 2
476 177
460 177
0 2 32 0 0 0 0 0 27 55 0 3
460 185
460 186
476 186
1 4 32 0 0 4224 0 15 27 0 0 3
460 135
460 204
470 204
3 0 33 0 0 4096 0 27 0 0 57 2
476 195
418 195
5 9 33 0 0 8320 0 18 28 0 0 3
418 229
418 180
284 180
14 4 19 0 0 0 0 28 18 0 0 2
278 243
367 243
2 3 34 0 0 4224 0 16 18 0 0 3
361 251
361 234
367 234
13 1 20 0 0 0 0 28 16 0 0 4
278 234
297 234
297 251
325 251
2 2 35 0 0 4224 0 17 18 0 0 2
363 225
367 225
12 1 21 0 0 0 0 28 17 0 0 2
278 225
327 225
11 1 22 0 0 0 0 28 18 0 0 2
278 216
367 216
0 4 36 0 0 8192 0 0 28 65 0 3
169 189
169 207
208 207
0 2 36 0 0 8192 0 0 28 66 0 3
169 180
169 189
214 189
1 1 36 0 0 4224 0 23 28 0 0 3
169 130
169 180
214 180
3 3 37 0 0 4224 0 24 28 0 0 2
98 198
214 198
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
