* C:\Users\gabriel\Desktop\SEMESTRE6\7.CE2Lab\projects\14-03.20-03\simulacoes\circuito1\circuit1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 26 16:41:44 2016



** Analysis setup **
.tran 0ns 10ms 0 20us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "circuit1.net"
.INC "circuit1.als"


.probe


.END
