CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
43032754 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 126 47 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
5 EWRED
-17 -26 18 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5130 0 0
2
42291.5 0
0
13 Logic Switch~
5 160 29 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
5 NSRED
-17 -26 18 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
391 0 0
2
42291.5 0
0
7 Ground~
168 140 366 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
42291.5 2
0
7 Pulser~
4 324 168 0 10 12
0 82 83 12 84 0 0 5 5 5
7
0
0 0 4640 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3421 0 0
2
42291.5 3
0
2 +V
167 919 266 0 1 3
0 20
0
0 0 54240 0
3 10V
29 -11 50 -3
2 V8
13 -11 27 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
42291.5 10
0
9 Inverter~
13 260 287 0 2 22
0 77 9
0
0 0 608 270
5 74F04
-18 -19 17 -11
4 U16A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
5572 0 0
2
42291.5 26
0
2 +V
167 79 164 0 1 3
0 39
0
0 0 54240 180
3 10V
6 -2 27 6
2 V1
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8901 0 0
2
42291.5 31
0
9 4-In AND~
219 468 244 0 5 22
0 53 56 52 54 43
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U11A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
7361 0 0
2
42291.5 32
0
9 Inverter~
13 388 218 0 2 22
0 55 53
0
0 0 608 0
5 74F04
-18 -30 17 -22
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
4747 0 0
2
42291.5 33
0
9 Inverter~
13 389 252 0 2 22
0 57 52
0
0 0 608 0
5 74F04
13 -17 48 -9
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
972 0 0
2
42291.5 34
0
9 Inverter~
13 387 340 0 2 22
0 51 46
0
0 0 608 0
5 74F04
13 -17 48 -9
4 U10A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3472 0 0
2
42291.5 35
0
9 Inverter~
13 388 302 0 2 22
0 49 47
0
0 0 608 0
5 74F04
-18 -30 17 -22
4 U10B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
9998 0 0
2
42291.5 36
0
9 4-In AND~
219 468 328 0 5 22
0 47 44 46 45 42
0
0 0 608 0
6 74LS21
-21 -28 21 -20
4 U11B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
3536 0 0
2
42291.5 37
0
9 Inverter~
13 354 359 0 2 22
0 48 45
0
0 0 608 0
5 74F04
13 -17 48 -9
4 U10C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
4597 0 0
2
42291.5 38
0
9 Inverter~
13 353 322 0 2 22
0 50 44
0
0 0 608 0
5 74F04
13 -17 48 -9
4 U10D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
3835 0 0
2
42291.5 39
0
9 2-In AND~
219 536 274 0 3 22
0 43 42 40
0
0 0 608 0
6 74LS08
-24 -36 18 -28
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3670 0 0
2
42291.5 40
0
6 74LS48
188 1022 79 0 14 29
0 55 56 57 54 95 96 65 64 63
62 61 60 59 97
0
0 0 4832 0
6 74LS48
-21 -76 21 -68
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
42291.5 41
0
9 Inverter~
13 929 148 0 2 22
0 56 66
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U7C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9323 0 0
2
42291.5 42
0
9 Inverter~
13 942 180 0 2 22
0 57 58
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U7B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
317 0 0
2
42291.5 43
0
9 Inverter~
13 694 146 0 2 22
0 49 67
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U7F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3108 0 0
2
42291.5 44
0
9 Inverter~
13 718 144 0 2 22
0 50 68
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U7E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
4299 0 0
2
42291.5 45
0
6 74LS48
188 814 78 0 14 29
0 49 50 51 48 98 99 75 74 73
72 71 70 69 100
0
0 0 4832 0
6 74LS48
-21 -76 21 -68
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
42291.5 46
0
10 4-In NAND~
219 617 94 0 5 22
0 54 58 66 55 76
0
0 0 608 180
6 74LS20
-21 -40 21 -32
3 U5A
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 1 0
1 U
7876 0 0
2
42291.5 47
0
9 CC 7-Seg~
183 88 244 0 12 19
10 69 70 71 72 73 74 75 2 2
0 1 1
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
5 DISP2
34 -4 69 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
6369 0 0
2
42291.5 48
0
9 CC 7-Seg~
183 193 243 0 16 19
10 59 60 61 62 63 64 65 2 2
1 1 0 1 1 0 1
0
0 0 21104 0
7 AMBERCC
-77 -28 -28 -20
5 DISP1
-70 -15 -35 -7
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
9172 0 0
2
42291.5 49
0
7 74LS160
124 145 139 0 14 29
0 39 39 76 39 101 102 103 104 78
105 49 50 51 48
0
0 0 4832 0
8 74LS160A
-25 -61 31 -53
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
7100 0 0
2
5.89727e-315 0
0
10 4-In NAND~
219 277 112 0 5 22
0 48 51 68 67 77
0
0 0 608 180
6 74LS20
-21 -40 21 -32
3 U5B
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
3820 0 0
2
5.89727e-315 5.26354e-315
0
14 Logic Display~
6 825 288 0 1 2
10 9
0
0 0 53872 0
6 100MEG
16 1 58 9
6 TMLONG
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89727e-315 5.30499e-315
0
2 +V
167 612 200 0 1 3
0 41
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
961 0 0
2
5.89727e-315 5.32571e-315
0
14 Logic Display~
6 749 287 0 1 2
10 10
0
0 0 53872 0
6 100MEG
16 1 58 9
7 TMSHORT
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89727e-315 5.34643e-315
0
10 2-In NAND~
219 264 38 0 3 22
0 8 7 80
0
0 0 608 0
4 7400
-15 -36 13 -28
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3409 0 0
2
5.89727e-315 5.3568e-315
0
9 2-In AND~
219 543 85 0 3 22
0 76 80 79
0
0 0 608 180
6 74LS08
-24 -36 18 -28
3 U9B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3951 0 0
2
5.89727e-315 5.36716e-315
0
9 2-In AND~
219 222 103 0 3 22
0 77 80 78
0
0 0 608 180
6 74LS08
-24 -36 18 -28
3 U9A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8885 0 0
2
5.89727e-315 5.37752e-315
0
7 74LS163
126 462 121 0 14 29
0 81 81 12 81 106 107 108 109 79
110 55 56 57 54
0
0 0 4832 0
8 74LS163A
-28 -62 28 -54
2 U2
-8 -52 6 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3780 0 0
2
5.89727e-315 5.38788e-315
0
5 7474~
219 612 292 0 6 22
0 41 41 40 78 111 10
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
9265 0 0
2
42291.5 50
0
2 +V
167 418 77 0 1 3
0 81
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
42291.5 51
0
121
8 0 2 0 0 8192 0 24 0 0 4 3
109 280
109 299
129 299
8 0 2 0 0 8192 0 25 0 0 3 3
214 279
214 299
242 299
1 9 2 0 0 8320 0 3 25 0 0 4
140 360
242 360
242 201
193 201
9 1 2 0 0 0 0 24 3 0 0 4
88 202
129 202
129 360
140 360
3 3 12 0 0 8320 0 4 34 0 0 4
348 159
385 159
385 112
430 112
2 1 7 0 0 0 0 31 1 0 0 2
240 47
138 47
1 1 8 0 0 0 0 31 2 0 0 2
240 29
172 29
4 0 39 0 0 4096 0 26 0 0 10 2
107 139
79 139
2 0 39 0 0 4096 0 26 0 0 10 2
113 121
79 121
1 1 39 0 0 8320 0 26 7 0 0 3
113 112
79 112
79 149
3 3 40 0 0 4224 0 16 35 0 0 2
557 274
588 274
2 1 9 0 0 8320 0 6 28 0 0 4
263 305
263 415
825 415
825 306
6 1 10 0 0 0 0 35 30 0 0 5
636 256
675 256
675 320
749 320
749 305
2 0 41 0 0 12416 0 35 0 0 15 4
588 256
575 256
575 220
612 220
1 1 41 0 0 0 0 29 35 0 0 2
612 209
612 229
5 2 42 0 0 8320 0 13 16 0 0 4
489 328
502 328
502 283
512 283
5 1 43 0 0 8320 0 8 16 0 0 4
489 244
502 244
502 265
512 265
2 2 44 0 0 12416 0 15 13 0 0 4
374 322
381 322
381 324
444 324
2 4 45 0 0 4224 0 14 13 0 0 4
375 359
429 359
429 342
444 342
2 3 46 0 0 12416 0 11 13 0 0 4
408 340
425 340
425 333
444 333
2 1 47 0 0 12416 0 12 13 0 0 4
409 302
425 302
425 315
444 315
0 1 48 0 0 4096 0 0 14 26 0 4
301 346
333 346
333 359
339 359
3 1 49 0 0 12288 0 0 12 26 0 4
301 311
316 311
316 302
373 302
2 1 50 0 0 4096 0 0 15 26 0 2
301 322
338 322
1 1 51 0 0 12288 0 0 11 26 0 4
301 336
316 336
316 340
372 340
1 0 1 0 0 4128 0 0 0 0 0 2
301 302
301 351
2 3 52 0 0 12416 0 10 8 0 0 4
410 252
425 252
425 249
444 249
2 1 53 0 0 12416 0 9 8 0 0 4
409 218
425 218
425 231
444 231
0 4 54 0 0 12288 0 0 8 33 0 6
301 262
333 262
333 275
429 275
429 258
444 258
3 1 55 0 0 12288 0 0 9 33 0 4
301 227
316 227
316 218
373 218
2 2 56 0 0 4224 0 0 8 33 0 4
301 238
381 238
381 240
444 240
1 1 57 0 0 4096 0 0 10 33 0 2
301 252
374 252
4 0 1 0 0 32 0 0 0 0 0 2
301 218
301 267
2 1 58 0 0 4224 0 19 0 0 48 2
945 198
945 248
13 0 59 0 0 4096 0 17 0 0 42 2
1054 97
1093 97
12 1 60 0 0 4096 0 17 0 0 42 2
1054 88
1093 88
11 2 61 0 0 4096 0 17 0 0 42 2
1054 79
1093 79
10 3 62 0 0 4096 0 17 0 0 42 2
1054 70
1093 70
9 4 63 0 0 4096 0 17 0 0 42 2
1054 61
1093 61
8 5 64 0 0 4096 0 17 0 0 42 2
1054 52
1093 52
7 6 65 0 0 4096 0 17 0 0 42 2
1054 43
1093 43
6 0 1 0 0 4256 0 0 0 0 0 2
1093 35
1093 106
0 3 55 0 0 4224 0 0 0 49 48 4
920 43
920 239
925 239
925 248
2 2 66 0 0 4224 0 18 0 0 48 2
932 166
932 248
0 0 54 0 0 4224 0 0 0 52 48 4
975 70
975 207
958 207
958 248
0 1 57 0 0 4224 0 0 19 51 0 2
945 61
945 162
0 1 56 0 0 0 0 0 18 50 0 2
932 52
932 130
5 0 1 0 0 32 0 0 0 0 0 2
915 248
969 248
3 1 55 0 0 0 0 0 17 53 0 2
910 43
990 43
2 2 56 0 0 0 0 0 17 53 0 2
910 52
990 52
1 3 57 0 0 0 0 0 17 53 0 2
910 61
990 61
0 4 54 0 0 0 0 0 17 53 0 2
910 70
990 70
4 0 1 0 0 32 0 0 0 0 0 2
910 26
910 75
2 3 67 0 0 4224 0 20 0 0 68 4
697 164
697 219
719 219
719 247
2 2 68 0 0 4224 0 21 0 0 68 4
721 162
721 208
728 208
728 247
0 1 49 0 0 4096 0 0 20 69 0 4
715 42
715 105
697 105
697 128
1 0 50 0 0 4096 0 21 0 0 70 2
721 126
721 51
13 0 69 0 0 4096 0 22 0 0 65 2
846 96
885 96
12 1 70 0 0 4096 0 22 0 0 65 2
846 87
885 87
11 2 71 0 0 4096 0 22 0 0 65 2
846 78
885 78
10 3 72 0 0 4096 0 22 0 0 65 2
846 69
885 69
9 4 73 0 0 4096 0 22 0 0 65 2
846 60
885 60
8 5 74 0 0 4096 0 22 0 0 65 2
846 51
885 51
7 6 75 0 0 4096 0 22 0 0 65 2
846 42
885 42
3 0 1 0 0 32 0 0 0 0 0 2
885 34
885 105
0 0 48 0 0 4224 0 0 0 72 68 2
748 69
748 247
1 0 51 0 0 4224 0 0 0 68 71 2
735 247
735 60
2 0 1 0 0 32 0 0 0 0 0 2
705 247
759 247
3 1 49 0 0 4224 0 0 22 73 0 2
700 42
782 42
2 2 50 0 0 4224 0 0 22 73 0 2
700 51
782 51
1 3 51 0 0 0 0 0 22 73 0 2
700 60
782 60
0 4 48 0 0 0 0 0 22 73 0 2
700 69
782 69
1 0 1 0 0 32 0 0 0 0 0 2
700 25
700 74
5 0 76 0 0 4096 0 23 0 0 111 2
590 94
568 94
1 0 54 0 0 0 0 23 0 0 79 2
641 107
671 107
4 3 55 0 0 0 0 23 0 0 79 2
641 80
671 80
2 1 58 0 0 0 0 23 0 0 79 2
641 98
671 98
3 2 66 0 0 0 0 23 0 0 79 2
641 89
671 89
5 0 1 0 0 32 0 0 0 0 0 2
671 64
671 120
1 0 59 0 0 4224 0 25 0 0 87 2
172 279
172 325
2 1 60 0 0 4224 0 25 0 0 87 2
178 279
178 325
3 2 61 0 0 4224 0 25 0 0 87 2
184 279
184 325
4 3 62 0 0 4224 0 25 0 0 87 2
190 279
190 325
5 4 63 0 0 4224 0 25 0 0 87 2
196 279
196 325
6 5 64 0 0 4224 0 25 0 0 87 2
202 279
202 325
7 6 65 0 0 4224 0 25 0 0 87 2
208 279
208 325
6 0 1 0 0 32 0 0 0 0 0 2
163 325
227 325
1 0 69 0 0 4224 0 24 0 0 95 2
67 280
67 326
2 1 70 0 0 4224 0 24 0 0 95 2
73 280
73 326
3 2 71 0 0 4224 0 24 0 0 95 2
79 280
79 326
4 3 72 0 0 4224 0 24 0 0 95 2
85 280
85 326
5 4 73 0 0 4224 0 24 0 0 95 2
91 280
91 326
6 5 74 0 0 4224 0 24 0 0 95 2
97 280
97 326
7 6 75 0 0 4224 0 24 0 0 95 2
103 280
103 326
3 0 1 0 0 32 0 0 0 0 0 2
58 326
122 326
1 0 48 0 0 0 0 27 0 0 100 2
301 125
334 125
2 1 51 0 0 0 0 27 0 0 100 2
301 116
334 116
3 2 68 0 0 0 0 27 0 0 100 2
301 107
334 107
4 3 67 0 0 0 0 27 0 0 100 2
301 98
334 98
2 0 1 0 0 32 0 0 0 0 0 2
334 82
334 138
0 1 77 0 0 12416 0 0 6 107 0 4
245 112
245 150
263 150
263 269
0 4 78 0 0 16512 0 0 35 104 0 6
183 103
183 70
48 70
48 387
612 387
612 304
9 3 79 0 0 8320 0 34 32 0 0 4
500 94
508 94
508 85
516 85
9 3 78 0 0 0 0 26 33 0 0 3
183 112
183 103
195 103
0 2 80 0 0 4224 0 0 32 106 0 4
308 38
587 38
587 76
561 76
3 2 80 0 0 0 0 31 33 0 0 6
291 38
309 38
309 71
257 71
257 94
240 94
5 1 77 0 0 0 0 27 33 0 0 2
250 112
240 112
1 0 81 0 0 4096 0 34 0 0 110 2
430 94
418 94
2 0 81 0 0 0 0 34 0 0 110 2
430 103
418 103
1 4 81 0 0 4224 0 36 34 0 0 3
418 86
418 121
424 121
1 3 76 0 0 12416 0 32 26 0 0 6
561 94
569 94
569 196
94 196
94 130
113 130
11 3 55 0 0 0 0 34 0 0 116 2
494 130
538 130
12 2 56 0 0 0 0 34 0 0 116 2
494 139
538 139
13 1 57 0 0 0 0 34 0 0 116 2
494 148
538 148
14 0 54 0 0 0 0 34 0 0 116 2
494 157
538 157
4 0 1 0 0 32 0 0 0 0 0 2
538 116
538 165
11 3 49 0 0 0 0 26 0 0 121 2
177 148
220 148
12 2 50 0 0 0 0 26 0 0 121 2
177 157
220 157
13 1 51 0 0 0 0 26 0 0 121 2
177 166
220 166
14 0 48 0 0 0 0 26 0 0 121 2
177 175
220 175
1 0 1 0 0 32 0 0 0 0 0 2
220 134
220 183
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
185 31 228 47
185 31 228 47
5 EWRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
188 13 231 29
188 13 231 29
5 NSRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 6
679 399 730 415
679 399 730 415
6 TMLONG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
676 304 735 320
676 304 735 320
7 TMSHORT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
