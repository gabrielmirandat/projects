CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 1 1
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
43032754 0
0
6 Title:
5 Name:
0
0
0
49
13 Logic Switch~
5 668 778 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21856 90
2 5V
14 -10 28 -2
3 V11
-10 -28 11 -20
3 FF3
10 0 31 8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8402 0 0
2
42269.8 0
0
13 Logic Switch~
5 630 779 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21856 90
2 5V
14 -10 28 -2
3 V10
-10 -28 11 -20
3 FF2
10 0 31 8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3751 0 0
2
42269.8 1
0
13 Logic Switch~
5 582 779 0 1 11
0 8
0
0 0 21856 90
2 0V
14 -10 28 -2
2 V9
-7 -28 7 -20
3 FF1
10 0 31 8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4292 0 0
2
42269.8 2
0
13 Logic Switch~
5 542 779 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21856 90
2 5V
11 -10 25 -2
2 V8
-7 -28 7 -20
2 PE
11 0 25 8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6118 0 0
2
42269.8 3
0
13 Logic Switch~
5 36 194 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
2 V7
-7 -28 7 -20
6 ENABLE
-20 -36 22 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
42269.8 4
0
13 Logic Switch~
5 31 305 0 1 11
0 16
0
0 0 22240 0
2 0V
-7 -18 7 -10
6 UPDOWN
-20 -28 22 -20
7 ENTRADA
-23 -39 26 -31
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6357 0 0
2
42269.8 5
0
13 Logic Switch~
5 493 778 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21856 90
2 5V
21 -10 35 -2
2 V1
-7 -28 7 -20
5 RESET
10 0 45 8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
319 0 0
2
42269.8 6
0
13 Logic Switch~
5 47 64 0 1 11
0 44
0
0 0 21856 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
12 CLOCK MANUAL
-41 -36 43 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3976 0 0
2
42269.8 7
0
8 2-In OR~
219 854 862 0 3 22
0 11 8 5
0
0 0 608 0
6 74LS32
-21 -36 21 -28
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
7634 0 0
2
5.89724e-315 0
0
8 2-In OR~
219 852 777 0 3 22
0 11 9 6
0
0 0 608 0
6 74LS32
-21 -37 21 -29
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
523 0 0
2
5.89724e-315 0
0
8 2-In OR~
219 851 696 0 3 22
0 11 10 7
0
0 0 608 0
6 74LS32
-21 -38 21 -30
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6748 0 0
2
5.89724e-315 0
0
9 2-In AND~
219 1198 655 0 3 22
0 5 12 2
0
0 0 2656 90
5 74F08
-18 -36 17 -28
3 U9C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
6901 0 0
2
5.89724e-315 0
0
9 2-In AND~
219 1135 655 0 3 22
0 6 12 3
0
0 0 2656 90
5 74F08
-18 -36 17 -28
3 U9B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
842 0 0
2
5.89724e-315 0
0
9 2-In AND~
219 1073 656 0 3 22
0 7 12 4
0
0 0 2656 90
5 74F08
-18 -36 17 -28
3 U9A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3277 0 0
2
5.89724e-315 0
0
10 3-In NAND~
219 720 385 0 4 22
0 13 12 10 21
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 7 0
1 U
4212 0 0
2
42269.8 8
0
10 3-In NAND~
219 718 268 0 4 22
0 13 12 9 14
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 7 0
1 U
4720 0 0
2
42269.8 9
0
10 3-In NAND~
219 718 57 0 4 22
0 13 12 8 15
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 7 0
1 U
5551 0 0
2
42269.8 10
0
9 Inverter~
13 603 47 0 2 22
0 11 13
0
0 0 608 0
5 74F04
-17 -30 18 -22
3 U8E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
6986 0 0
2
42269.8 11
0
9 2-In AND~
219 109 130 0 3 22
0 20 18 19
0
0 0 2656 0
5 74F08
-18 -36 17 -28
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8745 0 0
2
5.89724e-315 0
0
9 Inverter~
13 150 130 0 2 22
0 19 17
0
0 0 608 0
5 74F04
-17 -30 18 -22
3 U8D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
9592 0 0
2
42269.8 12
0
9 Inverter~
13 755 458 0 2 22
0 24 23
0
0 0 608 0
5 74F04
-18 -34 17 -26
3 U8C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
8748 0 0
2
42269.8 13
0
9 Inverter~
13 336 322 0 2 22
0 34 33
0
0 0 608 0
5 74F04
-18 -32 17 -24
3 U8B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
7168 0 0
2
5.89724e-315 5.26354e-315
0
9 Inverter~
13 338 261 0 2 22
0 39 38
0
0 0 608 0
5 74F04
-17 -30 18 -22
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
631 0 0
2
5.89724e-315 5.30499e-315
0
9 2-In XOR~
219 274 492 0 3 22
0 35 36 24
0
0 0 608 0
5 74F86
-18 -24 17 -16
3 U7B
-5 -35 16 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
9466 0 0
2
5.89724e-315 5.32571e-315
0
9 2-In XOR~
219 203 460 0 3 22
0 16 27 35
0
0 0 608 0
5 74F86
-18 -35 17 -27
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3266 0 0
2
5.89724e-315 5.34643e-315
0
9 2-In XOR~
219 210 405 0 3 22
0 16 27 32
0
0 0 608 0
5 74F86
-18 -37 17 -29
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
7693 0 0
2
5.89724e-315 5.3568e-315
0
9 2-In XOR~
219 208 339 0 3 22
0 16 27 34
0
0 0 608 0
5 74F86
-18 -35 17 -27
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3723 0 0
2
5.89724e-315 5.36716e-315
0
9 2-In XOR~
219 206 279 0 3 22
0 16 36 39
0
0 0 608 0
5 74F86
-18 -34 17 -26
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3440 0 0
2
5.89724e-315 5.37752e-315
0
9 2-In XOR~
219 205 223 0 3 22
0 16 36 37
0
0 0 608 0
5 74F86
-18 -35 17 -27
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
6263 0 0
2
5.89724e-315 5.38788e-315
0
9 3-In AND~
219 1147 296 0 4 22
0 27 26 25 41
0
0 0 608 0
5 74F11
-22 -36 13 -28
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
4900 0 0
2
5.89724e-315 5.39306e-315
0
9 2-In AND~
219 435 400 0 3 22
0 32 40 28
0
0 0 2656 0
5 74F08
-20 -37 15 -29
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
8783 0 0
2
5.89724e-315 5.39824e-315
0
9 2-In AND~
219 433 332 0 3 22
0 33 40 29
0
0 0 2656 0
5 74F08
-20 -37 15 -29
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3221 0 0
2
5.89724e-315 5.40342e-315
0
9 2-In AND~
219 430 236 0 3 22
0 38 25 30
0
0 0 2656 0
5 74F08
-17 -38 18 -30
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3215 0 0
2
5.89724e-315 5.4086e-315
0
9 2-In AND~
219 427 159 0 3 22
0 37 25 31
0
0 0 2656 0
5 74F08
-18 -36 17 -28
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7903 0 0
2
5.89724e-315 5.41378e-315
0
14 Logic Display~
6 936 413 0 1 2
10 25
0
0 0 53872 0
6 100MEG
0 -34 42 -26
2 Q3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7121 0 0
2
5.89724e-315 5.41896e-315
0
14 Logic Display~
6 910 411 0 1 2
10 40
0
0 0 53872 0
6 100MEG
-17 -32 25 -24
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
5.89724e-315 5.42414e-315
0
6 74112~
219 871 494 0 7 32
0 21 23 22 24 4 25 40
0
0 0 4704 0
5 74112
-41 -71 -6 -63
5 FFJK3
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
5996 0 0
2
5.89724e-315 5.42933e-315
0
6 74112~
219 876 337 0 7 32
0 14 29 22 28 3 26 36
0
0 0 4704 0
5 74112
-50 -67 -15 -59
5 FFJK2
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 6 0
1 U
7804 0 0
2
42269.8 14
0
6 74112~
219 876 195 0 7 32
0 15 31 22 30 2 42 27
0
0 0 4704 0
5 74112
4 -60 39 -52
5 FFJK1
-49 -71 -14 -63
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 6 0
1 U
5523 0 0
2
42269.8 15
0
14 Logic Display~
6 981 249 0 1 2
10 26
0
0 0 53872 0
6 100MEG
-54 -30 -12 -22
3 Q0b
-11 -30 10 -22
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
42269.8 16
0
14 Logic Display~
6 1027 102 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -32 45 -24
3 Q1b
26 -20 47 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
42269.8 17
0
14 Logic Display~
6 957 249 0 1 2
10 36
0
0 0 53872 0
6 100MEG
14 -22 56 -14
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
42269.8 18
0
14 Logic Display~
6 1005 102 0 1 2
10 27
0
0 0 53872 0
6 100MEG
-24 -35 18 -27
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
42269.8 19
0
14 Logic Display~
6 1200 142 0 1 2
10 41
0
0 0 54896 0
6 100MEG
10 -14 52 -6
1 S
20 -26 27 -18
6 ULTIMO
-21 -41 21 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
42269.8 20
0
14 Logic Display~
6 359 52 0 1 2
10 22
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 C
-13 -17 -6 -9
5 CLOCK
-9 -29 26 -21
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
42269.8 21
0
7 Pulser~
4 42 130 0 10 12
0 43 46 20 47 0 0 2 2 2
8
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7376 0 0
2
42269.8 22
0
2 +V
167 227 174 0 1 3
0 45
0
0 0 54240 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9156 0 0
2
42269.8 23
0
2 +V
167 227 26 0 1 3
0 43
0
0 0 54240 0
3 10V
9 -1 30 7
2 V1
11 -12 25 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5776 0 0
2
42269.8 24
0
5 7474~
219 227 139 0 6 22
0 43 44 17 45 48 22
0
0 0 864 0
4 7474
7 -73 35 -65
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
7207 0 0
2
42269.8 25
0
79
5 3 2 0 0 12432 0 39 12 0 0 5
876 207
876 210
1177 210
1177 631
1197 631
5 3 3 0 0 12416 0 38 13 0 0 4
876 349
876 370
1134 370
1134 631
5 3 4 0 0 8320 0 37 14 0 0 4
871 506
871 535
1072 535
1072 632
3 1 5 0 0 4224 0 9 12 0 0 3
887 862
1188 862
1188 676
3 1 6 0 0 4224 0 10 13 0 0 3
885 777
1125 777
1125 676
3 1 7 0 0 4224 0 11 14 0 0 3
884 696
1063 696
1063 677
2 0 8 0 0 8192 0 9 0 0 26 4
841 871
754 871
754 669
583 669
2 0 9 0 0 4096 0 10 0 0 21 4
839 786
714 786
714 745
631 745
2 0 10 0 0 4096 0 11 0 0 20 2
838 705
667 705
0 1 11 0 0 4096 0 0 9 11 0 3
799 766
799 853
841 853
0 1 11 0 0 0 0 0 10 12 0 3
799 687
799 768
839 768
1 0 11 0 0 4096 0 11 0 0 19 2
838 687
543 687
0 2 12 0 0 4096 0 0 12 14 0 3
1142 726
1206 726
1206 676
0 2 12 0 0 0 0 0 13 15 0 3
1081 726
1143 726
1143 676
2 0 12 0 0 8192 0 14 0 0 18 3
1081 677
1081 727
494 727
2 0 12 0 0 0 0 15 0 0 18 2
696 385
494 385
2 0 12 0 0 0 0 16 0 0 18 2
694 268
494 268
1 2 12 0 0 4224 0 7 17 0 0 3
494 765
494 57
694 57
1 1 11 0 0 8320 0 18 4 0 0 3
588 47
543 47
543 766
1 3 10 0 0 8320 0 1 15 0 0 4
669 765
667 765
667 394
696 394
1 3 9 0 0 4224 0 2 16 0 0 3
631 766
631 277
694 277
0 1 13 0 0 4096 0 0 15 23 0 3
637 259
637 376
696 376
0 1 13 0 0 4224 0 0 16 27 0 3
637 48
637 259
694 259
4 1 14 0 0 4224 0 16 38 0 0 4
745 268
875 268
875 274
876 274
1 4 15 0 0 8320 0 39 17 0 0 3
876 132
876 57
745 57
1 3 8 0 0 4224 0 3 17 0 0 3
583 766
583 66
694 66
2 1 13 0 0 0 0 18 17 0 0 4
624 47
637 47
637 48
694 48
1 0 16 0 0 4096 0 28 0 0 65 2
190 270
62 270
1 0 16 0 0 4096 0 27 0 0 31 2
192 330
61 330
1 0 16 0 0 4096 0 26 0 0 31 2
194 396
61 396
0 1 16 0 0 4224 0 0 25 65 0 3
61 305
61 451
187 451
2 3 17 0 0 12416 0 20 49 0 0 4
171 130
177 130
177 121
203 121
2 1 18 0 0 8320 0 19 5 0 0 4
85 139
73 139
73 194
48 194
3 1 19 0 0 4224 0 19 20 0 0 2
130 130
135 130
3 1 20 0 0 4224 0 46 19 0 0 2
66 121
85 121
4 1 21 0 0 4224 0 15 37 0 0 3
747 385
871 385
871 431
3 0 22 0 0 4096 0 39 0 0 70 2
846 168
807 168
2 2 23 0 0 4224 0 37 21 0 0 2
847 458
776 458
0 1 24 0 0 8192 0 0 21 47 0 3
618 476
618 458
740 458
0 3 25 0 0 8192 0 0 30 62 0 4
938 477
1100 477
1100 305
1123 305
0 2 26 0 0 4224 0 0 30 71 0 4
981 317
1077 317
1077 296
1123 296
0 1 27 0 0 8192 0 0 30 53 0 4
1004 159
1100 159
1100 287
1123 287
3 4 28 0 0 12416 0 31 38 0 0 4
456 400
532 400
532 319
852 319
2 3 29 0 0 4224 0 38 32 0 0 3
852 301
454 301
454 332
4 3 30 0 0 12416 0 39 33 0 0 4
852 177
762 177
762 236
451 236
2 3 31 0 0 4224 0 39 34 0 0 2
852 159
448 159
4 3 24 0 0 12416 0 37 24 0 0 4
847 476
618 476
618 492
307 492
3 1 32 0 0 12416 0 26 31 0 0 4
243 405
246 405
246 391
411 391
1 2 33 0 0 4224 0 32 22 0 0 4
409 323
372 323
372 322
357 322
3 1 34 0 0 12416 0 27 22 0 0 4
241 339
245 339
245 322
321 322
2 0 27 0 0 0 0 25 0 0 53 2
187 469
143 469
2 0 27 0 0 0 0 26 0 0 53 2
194 414
143 414
0 2 27 0 0 8320 0 0 27 74 0 5
1004 159
1004 617
143 617
143 348
192 348
3 1 35 0 0 8320 0 25 24 0 0 4
236 460
249 460
249 483
258 483
2 0 36 0 0 4096 0 24 0 0 60 2
258 501
169 501
3 1 37 0 0 4224 0 29 34 0 0 4
238 223
355 223
355 150
403 150
2 1 38 0 0 8320 0 23 33 0 0 4
359 261
374 261
374 227
406 227
3 1 39 0 0 12416 0 28 23 0 0 4
239 279
246 279
246 261
323 261
2 0 36 0 0 0 0 28 0 0 60 2
190 288
169 288
0 2 36 0 0 8320 0 0 29 73 0 5
957 299
957 596
169 596
169 232
189 232
2 0 25 0 0 0 0 33 0 0 62 4
406 245
390 245
390 279
380 279
0 2 25 0 0 8320 0 0 34 68 0 5
938 475
938 574
380 574
380 168
403 168
0 2 40 0 0 4096 0 0 31 64 0 4
401 407
416 407
416 409
411 409
0 2 40 0 0 8320 0 0 32 69 0 5
910 457
910 553
401 553
401 341
409 341
1 1 16 0 0 0 0 6 29 0 0 4
43 305
62 305
62 214
189 214
0 3 22 0 0 4096 0 0 37 70 0 3
807 305
807 467
841 467
4 1 41 0 0 8320 0 30 44 0 0 3
1168 296
1200 296
1200 160
1 6 25 0 0 0 0 35 37 0 0 4
936 431
938 431
938 476
901 476
7 1 40 0 0 0 0 37 36 0 0 3
895 458
910 458
910 429
0 3 22 0 0 4224 0 0 38 75 0 4
358 103
807 103
807 310
846 310
6 1 26 0 0 0 0 38 40 0 0 3
906 319
981 319
981 267
6 1 42 0 0 4224 0 39 41 0 0 3
906 177
1027 177
1027 120
7 1 36 0 0 0 0 38 42 0 0 3
900 301
957 301
957 267
7 1 27 0 0 0 0 39 43 0 0 4
900 159
1006 159
1006 120
1005 120
6 1 22 0 0 0 0 49 45 0 0 3
251 103
359 103
359 70
0 1 43 0 0 4224 0 0 46 79 0 4
227 39
8 39
8 121
18 121
1 2 44 0 0 4224 0 8 49 0 0 4
59 64
188 64
188 103
203 103
4 1 45 0 0 4224 0 49 47 0 0 2
227 151
227 159
1 1 43 0 0 0 0 48 49 0 0 2
227 35
227 76
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
