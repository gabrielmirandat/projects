CircuitMaker Text
5.6
Probes: 70
L4_2
AC Analysis
15 887 752 16711935
L4_2
DC Sweep
15 887 752 16711935
L4_2
Fourier Analysis
15 887 752 16711935
V8_1
AC Analysis
14 728 752 16776960
V8_1
DC Sweep
14 728 752 16776960
V8_1
Fourier Analysis
14 728 752 16776960
L3_2
AC Analysis
13 878 531 65535
L3_2
DC Sweep
13 878 531 65535
L3_2
Fourier Analysis
13 878 531 65535
V7_1
AC Analysis
12 738 531 65280
V7_1
DC Sweep
12 738 531 65280
V7_1
Fourier Analysis
12 738 531 65280
R6_2
AC Analysis
11 866 338 255
R6_2
DC Sweep
11 866 338 255
R6_2
Fourier Analysis
11 866 338 255
V4_1
AC Analysis
10 730 338 16711680
V4_1
DC Sweep
10 730 338 16711680
V4_1
Fourier Analysis
10 730 338 16711680
R5_2
AC Analysis
9 882 90 43690
R5_2
DC Sweep
9 882 90 43690
R5_2
Fourier Analysis
9 882 90 43690
V3_1
AC Analysis
8 739 90 32768
V3_1
DC Sweep
8 739 90 32768
V3_1
Fourier Analysis
8 739 90 32768
C4_2
AC Analysis
7 363 750 7829503
C4_2
DC Sweep
7 363 750 7829503
C4_2
Fourier Analysis
7 363 750 7829503
V6_1
AC Analysis
6 225 750 16742263
V6_1
DC Sweep
6 225 750 16742263
V6_1
Fourier Analysis
6 225 750 16742263
C3_2
AC Analysis
5 362 534 33023
C3_2
DC Sweep
5 362 534 33023
C3_2
Fourier Analysis
5 362 534 33023
V5_1
AC Analysis
4 220 534 11184640
V5_1
DC Sweep
4 220 534 11184640
V5_1
Fourier Analysis
4 220 534 11184640
C2_2
AC Analysis
3 361 330 16711935
C2_2
DC Sweep
3 361 330 16711935
C2_2
Fourier Analysis
3 361 330 16711935
V1_1
AC Analysis
2 236 330 16776960
V1_1
DC Sweep
2 236 330 16776960
V1_1
Fourier Analysis
2 236 330 16776960
C1_2
AC Analysis
1 386 85 65535
C1_2
DC Sweep
1 386 85 65535
C1_2
Fourier Analysis
1 386 85 65535
V2_1
AC Analysis
0 240 85 65280
V2_1
DC Sweep
0 240 85 65280
V2_1
Fourier Analysis
0 240 85 65280
V2_1
Operating Point
0 251 89 65280
C1_2
Operating Point
1 347 85 65535
V1_1
Operating Point
2 362 232 16776960
R2_2
Operating Point
3 463 230 16711935
V5_1
Operating Point
4 253 370 11184640
C3_2
Operating Point
5 354 373 33023
V6_1
Operating Point
6 348 517 16742263
C4_2
Operating Point
7 446 517 7829503
V3_1
Operating Point
8 713 93 32768
L1_2
Operating Point
9 842 92 43690
V4_1
Operating Point
10 844 229 16711680
R6_2
Operating Point
11 945 228 255
V7_1
Operating Point
12 726 373 65280
L3_2
Operating Point
13 820 374 65535
V8_1
Operating Point
14 823 515 16776960
L4_2
Operating Point
15 957 514 16711935
V4_1
Transient Analysis
10 841 230 16711680
R6_2
Transient Analysis
11 970 228 255
V7_1
Transient Analysis
12 730 369 65280
L3_2
Transient Analysis
13 835 371 65535
V8_1
Transient Analysis
14 831 513 16776960
L4_2
Transient Analysis
15 951 513 16711935
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 1 1
20 Package,Description,
93 C:\Users\Marina\Documents\4� semestre\Sistemas digitais 1\Laborat�rio\CircuitMakerfim\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
1083703314 0
0
6 Title:
5 Name:
0
0
0
48
11 Signal Gen~
195 699 570 0 64 64
0 4 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1229080480 0 1073846682
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 18
20
0 795770 0 2.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V8
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 2.025 795.8k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
5.8973e-315 5.34643e-315
0
5 SAVE-
218 957 515 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 P
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
391 0 0
2
5.8973e-315 5.32571e-315
0
5 SAVE-
218 815 516 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 O
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3124 0 0
2
5.8973e-315 5.30499e-315
0
7 Ground~
168 880 644 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
5.8973e-315 5.26354e-315
0
9 Inductor~
219 882 516 0 2 5
0 4 3
0
0 0 832 0
3 1mH
-11 -17 10 -9
2 L4
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.8973e-315 0
0
7 Ground~
168 773 213 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
5.8973e-315 5.3568e-315
0
9 Inductor~
219 771 91 0 2 5
0 6 5
0
0 0 832 0
3 1mH
-11 -17 10 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.8973e-315 5.32571e-315
0
11 Signal Gen~
195 592 139 0 64 64
0 6 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112047697 -1073636966 1073846682
0 814313567 814313567 1008953853 1017343536 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 254
20
0 50.1253 -2.025 2.025 0 1e-09 1e-09 0.009974 0.01995 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V3
-7 -40 7 -32
0
0
55 %D %1 %2 DC 0 PULSE(-2.025 2.025 0 1n 1n 9.974m 19.95m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.8973e-315 5.30499e-315
0
5 SAVE-
218 710 91 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 I
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4747 0 0
2
5.8973e-315 5.26354e-315
0
5 SAVE-
218 853 91 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 J
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
972 0 0
2
5.8973e-315 0
0
11 Signal Gen~
195 602 426 0 19 64
0 8 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1209756800 0 1073846682
20
0 159154 0 2.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V7
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 2.025 159.2k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.8973e-315 5.34643e-315
0
5 SAVE-
218 856 372 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 N
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9998 0 0
2
5.8973e-315 5.32571e-315
0
5 SAVE-
218 727 372 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 M
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3536 0 0
2
5.8973e-315 5.30499e-315
0
7 Ground~
168 783 497 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.8973e-315 5.26354e-315
0
9 Inductor~
219 785 372 0 2 5
0 8 7
0
0 0 832 0
3 1mH
-11 -17 10 -9
2 L3
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.8973e-315 0
0
11 Signal Gen~
195 216 570 0 64 64
0 10 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1173925274 0 1073846682
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 262
20
0 7957.7 0 2.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V6
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 2.025 7.958k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.8973e-315 5.34643e-315
0
5 SAVE-
218 473 516 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 H
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5616 0 0
2
5.8973e-315 5.32571e-315
0
5 SAVE-
218 335 516 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 G
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9323 0 0
2
5.8973e-315 5.30499e-315
0
10 Capacitor~
219 523 567 0 2 5
0 2 9
0
0 0 832 90
5 0.1uF
10 3 45 11
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
317 0 0
2
5.8973e-315 5.26354e-315
0
7 Ground~
168 394 644 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
5.8973e-315 0
0
7 Ground~
168 297 216 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4299 0 0
2
5.8973e-315 5.3568e-315
0
10 Capacitor~
219 426 139 0 2 5
0 2 11
0
0 0 832 90
5 0.1uF
10 3 45 11
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9672 0 0
2
5.8973e-315 5.32571e-315
0
11 Signal Gen~
195 116 142 0 64 64
0 12 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1140498534 -1073636966 1073846682
0 814313567 814313567 981642693 990035596 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 62
20
0 501.253 -2.025 2.025 0 1e-09 1e-09 0.000997 0.001995 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V2
-7 -40 7 -32
0
0
53 %D %1 %2 DC 0 PULSE(-2.025 2.025 0 1n 1n 997u 1.995m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
5.8973e-315 5.30499e-315
0
5 SAVE-
218 230 88 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
6369 0 0
2
5.8973e-315 5.26354e-315
0
5 SAVE-
218 376 88 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9172 0 0
2
5.8973e-315 0
0
11 Signal Gen~
195 113 426 0 64 64
0 14 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1153888584 0 1073846682
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 1591.54 0 2.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V5
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 2.025 1.592k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
5.8973e-315 5.34643e-315
0
5 SAVE-
218 362 372 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 E
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3820 0 0
2
5.8973e-315 5.32571e-315
0
5 SAVE-
218 220 372 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 F
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7678 0 0
2
5.8973e-315 5.30499e-315
0
10 Capacitor~
219 423 423 0 2 5
0 2 13
0
0 0 832 90
5 0.1uF
10 3 45 11
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
961 0 0
2
5.8973e-315 5.26354e-315
0
7 Ground~
168 294 497 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
5.8973e-315 0
0
7 Ground~
168 394 357 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
5.8973e-315 0
0
5 SAVE-
218 453 231 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 D
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3951 0 0
2
5.8973e-315 5.34643e-315
0
5 SAVE-
218 328 231 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
8885 0 0
2
5.8973e-315 5.32571e-315
0
11 Signal Gen~
195 213 285 0 64 64
0 16 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1134503789 0 1073846682
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 262
20
0 318.308 0 2.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 2.025 318.3 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3780 0 0
2
5.8973e-315 5.30499e-315
0
10 Capacitor~
219 523 282 0 2 5
0 2 15
0
0 0 832 90
5 0.1uF
10 3 45 11
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9265 0 0
2
5.8973e-315 5.26354e-315
0
11 Signal Gen~
195 706 283 0 64 64
0 18 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1190702490 0 1073846682
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 31830.8 0 2.025 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -2.02/2.02V
-38 -30 39 -22
2 V4
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 2.025 31.83k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
5.8973e-315 5.3568e-315
0
5 SAVE-
218 958 229 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 L
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9424 0 0
2
5.8973e-315 5.34643e-315
0
5 SAVE-
218 822 229 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 K
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
9968 0 0
2
5.8973e-315 5.32571e-315
0
9 Inductor~
219 889 229 0 2 5
0 18 17
0
0 0 832 0
3 1mH
-11 -17 10 -9
2 L2
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.8973e-315 5.30499e-315
0
7 Ground~
168 887 358 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8464 0 0
2
5.8973e-315 5.26354e-315
0
9 Resistor~
219 1016 567 0 3 5
0 2 3 -1
0
0 0 864 90
2 1k
15 0 29 8
2 R8
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7168 0 0
2
5.8973e-315 5.3568e-315
0
9 Resistor~
219 902 139 0 3 5
0 2 5 -1
0
0 0 864 90
2 1k
15 0 29 8
2 R5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3171 0 0
2
5.8973e-315 5.34643e-315
0
9 Resistor~
219 919 423 0 3 5
0 2 7 -1
0
0 0 864 90
2 1k
14 0 28 8
2 R7
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
4139 0 0
2
5.8973e-315 5.3568e-315
0
9 Resistor~
219 397 516 0 2 5
0 10 9
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
6435 0 0
2
5.8973e-315 5.3568e-315
0
9 Resistor~
219 300 88 0 2 5
0 12 11
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
5283 0 0
2
5.8973e-315 5.34643e-315
0
9 Resistor~
219 297 372 0 2 5
0 14 13
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
6874 0 0
2
5.8973e-315 5.3568e-315
0
9 Resistor~
219 397 231 0 2 5
0 16 15
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
5305 0 0
2
5.8973e-315 0
0
9 Resistor~
219 1023 280 0 3 5
0 2 17 -1
0
0 0 864 90
2 1k
15 0 29 8
2 R6
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
34 0 0
2
5.8973e-315 0
0
32
0 2 2 0 0 4096 0 0 1 3 0 4
880 616
758 616
758 575
730 575
2 2 3 0 0 4224 0 5 41 0 0 3
900 516
1016 516
1016 549
1 1 2 0 0 8192 0 41 4 0 0 4
1016 585
1016 616
880 616
880 638
1 1 4 0 0 12416 0 1 5 0 0 4
730 565
758 565
758 516
864 516
0 2 2 0 0 0 0 0 8 7 0 4
773 185
651 185
651 144
623 144
2 2 5 0 0 4224 0 7 42 0 0 3
789 91
902 91
902 121
1 1 2 0 0 0 0 42 6 0 0 4
902 157
902 185
773 185
773 207
1 1 6 0 0 12416 0 8 7 0 0 4
623 134
651 134
651 91
753 91
0 2 2 0 0 0 0 0 11 11 0 4
783 472
661 472
661 431
633 431
2 2 7 0 0 4224 0 15 43 0 0 3
803 372
919 372
919 405
1 1 2 0 0 0 0 43 14 0 0 4
919 441
919 472
783 472
783 491
1 1 8 0 0 12416 0 11 15 0 0 4
633 421
661 421
661 372
767 372
0 1 2 0 0 0 0 0 20 15 0 2
394 616
394 638
2 2 9 0 0 4224 0 44 19 0 0 3
415 516
523 516
523 558
2 1 2 0 0 12416 0 16 19 0 0 5
247 575
272 575
272 616
523 616
523 576
1 1 10 0 0 12416 0 16 44 0 0 4
247 565
272 565
272 516
379 516
0 1 2 0 0 0 0 0 21 19 0 2
297 188
297 210
2 2 11 0 0 4224 0 45 22 0 0 3
318 88
426 88
426 130
2 1 2 0 0 0 0 23 22 0 0 5
147 147
175 147
175 188
426 188
426 148
1 1 12 0 0 12416 0 23 45 0 0 4
147 137
175 137
175 88
282 88
0 1 2 0 0 0 0 0 30 23 0 2
294 472
294 491
2 2 13 0 0 4224 0 46 29 0 0 3
315 372
423 372
423 414
2 1 2 0 0 0 0 26 29 0 0 5
144 431
172 431
172 472
423 472
423 432
1 1 14 0 0 12416 0 26 46 0 0 4
144 421
172 421
172 372
279 372
0 1 2 0 0 0 0 0 31 27 0 2
394 331
394 351
2 2 15 0 0 4224 0 47 35 0 0 3
415 231
523 231
523 273
2 1 2 0 0 0 0 34 35 0 0 5
244 290
272 290
272 331
523 331
523 291
1 1 16 0 0 12416 0 34 47 0 0 4
244 280
272 280
272 231
379 231
0 2 2 0 0 0 0 0 36 31 0 4
887 329
765 329
765 288
737 288
2 2 17 0 0 4224 0 39 48 0 0 3
907 229
1023 229
1023 262
1 1 2 0 0 0 0 48 40 0 0 4
1023 298
1023 329
887 329
887 352
1 1 18 0 0 12416 0 36 39 0 0 4
737 278
765 278
765 229
871 229
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
