CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 210 5 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
176 393 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
10
5 SCOPE
12 760 267 0 1 11
0 2
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5130 0 0
2
42186.3 0
0
14 Logic Display~
6 785 218 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
391 0 0
2
42186.3 0
0
9 Inverter~
13 688 278 0 2 22
0 3 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3124 0 0
2
42186.3 0
0
12 Hex Display~
7 397 439 0 16 19
10 7 6 5 4 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3421 0 0
2
42186.3 0
0
5 4012~
219 569 301 0 5 22
0 4 5 9 8 3
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 2 0
1 U
8157 0 0
2
42186.3 0
0
9 Inverter~
13 455 342 0 2 22
0 7 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5572 0 0
2
42186.3 0
0
9 Inverter~
13 456 317 0 2 22
0 6 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8901 0 0
2
42186.3 0
0
2 +V
167 289 204 0 1 3
0 10
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
42186.3 0
0
7 74LS163
126 340 288 0 14 29
0 10 10 11 10 12 13 14 15 3
16 4 5 6 7
0
0 0 4848 0
8 74LS163A
-28 -51 28 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
4747 0 0
2
42186.3 0
0
7 Pulser~
4 149 290 0 10 12
0 17 18 11 19 0 0 10 10 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
972 0 0
2
42186.3 0
0
18
1 0 2 0 0 4096 0 1 0 0 2 2
760 279
760 278
2 1 2 0 0 4224 0 3 2 0 0 3
709 278
785 278
785 236
0 1 3 0 0 4096 0 0 3 8 0 2
596 278
673 278
0 4 4 0 0 4096 0 0 4 9 0 6
402 297
402 402
371 402
371 476
388 476
388 463
0 3 5 0 0 4096 0 0 4 10 0 6
411 306
411 407
376 407
376 471
394 471
394 463
0 2 6 0 0 4224 0 0 4 13 0 4
420 315
420 476
400 476
400 463
0 1 7 0 0 8320 0 0 4 14 0 5
432 342
419 342
419 471
406 471
406 463
5 9 3 0 0 8320 0 5 9 0 0 3
596 301
596 261
378 261
11 1 4 0 0 4224 0 9 5 0 0 4
372 297
537 297
537 288
545 288
12 2 5 0 0 12416 0 9 5 0 0 4
372 306
437 306
437 297
545 297
2 4 8 0 0 4224 0 6 5 0 0 4
476 342
532 342
532 315
545 315
2 3 9 0 0 4224 0 7 5 0 0 4
477 317
537 317
537 306
545 306
13 1 6 0 0 0 0 9 7 0 0 4
372 315
433 315
433 317
441 317
14 1 7 0 0 0 0 9 6 0 0 4
372 324
432 324
432 342
440 342
0 4 10 0 0 4096 0 0 9 16 0 3
289 270
289 288
302 288
0 2 10 0 0 8192 0 0 9 17 0 3
289 261
289 270
308 270
1 1 10 0 0 4224 0 8 9 0 0 3
289 213
289 261
308 261
3 3 11 0 0 4224 0 10 9 0 0 4
173 281
294 281
294 279
308 279
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
