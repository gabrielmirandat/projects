CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
353 178 1368 715
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
521 274 634 371
9478322 0
0
6 Title:
5 Name:
0
0
0
7
9 V Source~
197 543 239 0 1 5
0 0
0
0 0 17248 0
2 4V
16 0 30 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
5130 0 0
2
42282 0
0
9 V Source~
197 96 206 0 1 5
0 0
0
0 0 17248 0
2 6V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
391 0 0
2
42282 0
0
9 Resistor~
219 721 209 0 1 5
0 0
0
0 0 864 90
4 2.2k
1 0 29 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66071556
82 0 0 0 1 0 0 0
1 R
3124 0 0
2
42282 0
0
9 Resistor~
219 542 177 0 1 5
0 0
0
0 0 864 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66070708
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
42282 0
0
9 Resistor~
219 402 128 0 1 5
0 0
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66069844
82 0 0 0 1 0 0 0
1 R
8157 0 0
2
42282 0
0
9 Resistor~
219 288 206 0 1 5
0 0
0
0 0 864 90
4 4.7k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66069048
82 0 0 0 1 0 0 0
1 R
5572 0 0
2
42282 0
0
9 Resistor~
219 188 127 0 1 5
0 0
0
0 0 864 0
3 100
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66072404
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
42282 0
0
9
0 2 0 0 0 0 0 0 2 2 0 3
289 293
96 293
96 227
0 1 0 0 0 0 0 0 6 3 0 3
543 293
288 293
288 224
2 1 0 0 0 0 0 1 3 0 0 4
543 260
543 293
721 293
721 227
1 1 0 0 0 0 0 4 1 0 0 3
542 195
543 195
543 218
2 0 0 0 0 0 0 4 0 0 6 2
542 159
542 128
1 2 0 0 0 0 0 5 3 0 0 3
420 128
721 128
721 191
2 0 0 0 0 0 0 6 0 0 8 2
288 188
288 128
2 2 0 0 0 0 0 7 5 0 0 3
206 127
206 128
384 128
1 1 0 0 0 0 0 2 7 0 0 3
96 185
96 127
170 127
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
