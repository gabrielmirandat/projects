CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.433121 0.500000
344 175 1532 447
1083744434 0
0
6 Title:
5 Name:
0
0
0
9
7 Ground~
168 528 396 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
42282 0
0
8 Battery~
219 500 321 0 2 5
0 3 2
0
0 0 880 0
4 3.5V
9 -2 37 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
391 0 0
2
42282 0
0
9 Resistor~
219 889 166 0 3 5
0 2 4 -1
0
0 0 880 90
2 2k
8 0 22 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66204440
82 0 0 0 1 0 0 0
1 R
3124 0 0
2
42282 0
0
9 Resistor~
219 719 163 0 3 5
0 2 4 -1
0
0 0 880 90
2 2k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66203576
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
42282 0
0
9 Resistor~
219 615 127 0 2 5
0 4 5
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66202696
82 0 0 0 1 0 0 0
1 R
8157 0 0
2
42282 0
0
9 Resistor~
219 499 165 0 2 5
0 3 5
0
0 0 880 90
2 2k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66201868
82 0 0 0 1 0 0 0
1 R
5572 0 0
2
42282 0
0
9 Resistor~
219 405 126 0 2 5
0 6 5
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66201092
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
42282 0
0
9 Resistor~
219 291 166 0 2 5
0 3 6
0
0 0 880 90
2 2k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66200316
82 0 0 0 1 0 0 0
1 R
7361 0 0
2
42282 0
0
9 Resistor~
219 138 165 0 3 5
0 2 6 -1
0
0 0 880 90
2 2k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66212264
82 0 0 0 1 0 0 0
1 R
4747 0 0
2
42282 0
0
13
0 0 3 0 0 4096 0 0 0 3 0 3
500 292
634 292
634 258
1 0 2 0 0 12288 0 4 0 0 12 4
719 181
719 247
683 247
683 353
0 1 3 0 0 0 0 0 6 4 0 3
500 292
499 292
499 183
1 1 3 0 0 8320 0 2 8 0 0 6
500 308
500 292
349 292
349 267
291 267
291 184
1 0 2 0 0 0 0 1 0 0 12 2
528 390
528 353
2 0 4 0 0 4096 0 4 0 0 9 2
719 145
719 127
2 0 5 0 0 4096 0 6 0 0 10 2
499 147
499 127
2 0 6 0 0 4096 0 8 0 0 11 2
291 148
291 126
1 2 4 0 0 4224 0 5 3 0 0 3
633 127
889 127
889 148
2 2 5 0 0 8320 0 7 5 0 0 3
423 126
423 127
597 127
2 1 6 0 0 8320 0 9 7 0 0 3
138 147
138 126
387 126
0 1 2 0 0 4224 0 0 3 13 0 3
499 353
889 353
889 184
1 2 2 0 0 0 0 9 2 0 0 4
138 183
138 353
500 353
500 332
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
521 276 540 292
521 276 540 292
2 v4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
326 337 345 353
326 337 345 353
2 v0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
672 111 691 127
672 111 691 127
2 v3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
450 111 469 127
450 111 469 127
2 v2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
138 110 157 126
138 110 157 126
2 v1
0
17 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
