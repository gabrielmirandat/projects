CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
259 95 1274 632
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
427 191 540 288
43024402 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 42 272 0 1 11
0 7
0
0 0 22368 0
2 0V
-6 -16 8 -8
1 M
-3 -26 4 -18
5 MOEDA
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89721e-315 0
0
13 Logic Switch~
5 244 521 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
2 V1
-7 -28 7 -20
5 RESET
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89721e-315 5.26354e-315
0
13 Logic Switch~
5 92 103 0 1 11
0 17
0
0 0 21856 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
12 CLOCK MANUAL
-41 -36 43 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89721e-315 5.30499e-315
0
8 2-In OR~
219 343 401 0 3 22
0 7 4 6
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3421 0 0
2
5.89721e-315 5.32571e-315
0
8 2-In OR~
219 346 272 0 3 22
0 7 5 8
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8157 0 0
2
5.89721e-315 5.34643e-315
0
6 74112~
219 602 474 0 7 32
0 14 3 10 6 13 2 5
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U5B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 6 0
1 U
5572 0 0
2
5.89721e-315 5.3568e-315
0
6 74112~
219 602 227 0 7 32
0 9 8 10 9 13 3 4
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 6 0
1 U
8901 0 0
2
5.89721e-315 5.36716e-315
0
9 2-In AND~
219 832 360 0 3 22
0 4 2 11
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7361 0 0
2
5.89721e-315 5.37752e-315
0
9 2-In AND~
219 831 191 0 3 22
0 4 5 12
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4747 0 0
2
5.89721e-315 5.38788e-315
0
14 Logic Display~
6 684 386 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Q0b
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89721e-315 5.39306e-315
0
14 Logic Display~
6 688 142 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Q1b
-11 -20 10 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89721e-315 5.39824e-315
0
14 Logic Display~
6 652 388 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89721e-315 5.40342e-315
0
14 Logic Display~
6 651 143 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.89721e-315 5.4086e-315
0
2 +V
167 602 348 0 1 3
0 14
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4597 0 0
2
5.89721e-315 5.41378e-315
0
2 +V
167 602 102 0 1 3
0 9
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
5.89721e-315 5.41896e-315
0
14 Logic Display~
6 971 283 0 1 2
10 11
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 E
20 -26 27 -18
4 ERRO
-14 -41 14 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89721e-315 5.42414e-315
0
14 Logic Display~
6 972 136 0 1 2
10 12
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 R
20 -26 27 -18
7 RETORNO
-24 -41 25 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.89721e-315 5.42933e-315
0
14 Logic Display~
6 359 52 0 1 2
10 10
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
5 CLOCK
-18 -41 17 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89721e-315 5.43192e-315
0
7 Pulser~
4 82 157 0 10 12
0 16 19 15 20 0 0 2 2 2
7
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
317 0 0
2
5.89721e-315 5.43451e-315
0
2 +V
167 228 215 0 1 3
0 18
0
0 0 54240 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
5.89721e-315 5.4371e-315
0
2 +V
167 227 31 0 1 3
0 16
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
5.89721e-315 5.43969e-315
0
5 7474~
219 227 139 0 6 22
0 16 17 15 18 21 10
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9672 0 0
2
5.89721e-315 5.44228e-315
0
30
0 2 2 0 0 4224 0 0 8 2 0 4
684 456
795 456
795 369
808 369
6 1 2 0 0 0 0 6 10 0 0 3
632 456
684 456
684 404
0 2 3 0 0 12416 0 0 6 4 0 5
688 209
688 308
565 308
565 438
578 438
6 1 3 0 0 0 0 7 11 0 0 3
632 209
688 209
688 160
1 0 4 0 0 4096 0 8 0 0 8 2
808 351
720 351
0 2 5 0 0 8192 0 0 9 11 0 4
652 557
775 557
775 200
807 200
0 1 4 0 0 8192 0 0 9 8 0 4
720 275
784 275
784 182
807 182
0 2 4 0 0 16512 0 0 4 20 0 7
651 191
651 275
720 275
720 581
150 581
150 410
330 410
4 3 6 0 0 4224 0 6 4 0 0 4
578 456
458 456
458 401
376 401
0 1 7 0 0 8192 0 0 4 13 0 3
151 272
151 392
330 392
0 2 5 0 0 8320 0 0 5 19 0 5
652 438
652 557
187 557
187 281
333 281
2 3 8 0 0 4224 0 7 5 0 0 4
578 191
460 191
460 272
379 272
1 1 7 0 0 12416 0 1 5 0 0 4
54 272
152 272
152 263
333 263
0 4 9 0 0 4224 0 0 7 24 0 4
602 132
521 132
521 209
578 209
0 3 10 0 0 4224 0 0 6 16 0 3
544 200
544 447
572 447
0 3 10 0 0 0 0 0 7 25 0 4
359 103
544 103
544 200
572 200
3 1 11 0 0 4224 0 8 16 0 0 3
853 360
971 360
971 301
3 1 12 0 0 4224 0 9 17 0 0 3
852 191
972 191
972 154
7 1 5 0 0 0 0 6 12 0 0 3
626 438
652 438
652 406
7 1 4 0 0 0 0 7 13 0 0 3
626 191
651 191
651 161
5 0 13 0 0 12288 0 7 0 0 22 4
602 239
602 293
523 293
523 521
1 5 13 0 0 4224 0 2 6 0 0 3
256 521
602 521
602 486
1 1 14 0 0 4224 0 14 6 0 0 2
602 357
602 411
1 1 9 0 0 0 0 15 7 0 0 2
602 111
602 164
6 1 10 0 0 0 0 22 18 0 0 3
251 103
359 103
359 70
3 3 15 0 0 12416 0 19 22 0 0 4
106 148
151 148
151 121
203 121
0 1 16 0 0 4224 0 0 19 30 0 4
227 48
28 48
28 148
58 148
1 2 17 0 0 4224 0 3 22 0 0 2
104 103
203 103
4 1 18 0 0 4224 0 22 20 0 0 3
227 151
227 200
228 200
1 1 16 0 0 0 0 21 22 0 0 2
227 40
227 76
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
