* C:\Users\Marina\Desktop\EXP6C.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 27 13:12:33 2015



** Analysis setup **
.tran 1ns 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EXP6C.net"
.INC "EXP6C.als"


.probe


.END
