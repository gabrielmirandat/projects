* C:\Users\gabriel\Dropbox\SEMESTRE6\7.CE2Lab\projects\proj4\passa-baixas\passa_baixas.sch

* Schematics Version 9.1 - Web Update 1
* Thu Apr 28 13:14:12 2016



** Analysis setup **
.tran 0ns 10ms 0 20us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "passa_baixas.net"
.INC "passa_baixas.als"


.probe


.END
