CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 C:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 92 210 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
733 0 0
2
42183 0
0
13 Logic Switch~
5 96 169 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9115 0 0
2
42183 0
0
13 Logic Switch~
5 97 123 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4192 0 0
2
42183 0
0
14 Logic Display~
6 482 95 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4509 0 0
2
42183 0
0
14 Logic Display~
6 443 96 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9887 0 0
2
42183 0
0
10 2-In NAND~
219 351 205 0 3 22
0 2 4 3
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6657 0 0
2
42183 0
0
10 2-In NAND~
219 353 139 0 3 22
0 5 3 2
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6962 0 0
2
42183 0
0
10 2-In NAND~
219 228 209 0 3 22
0 6 7 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3881 0 0
2
42183 0
0
10 2-In NAND~
219 225 133 0 3 22
0 8 6 5
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3536 0 0
2
42183 0
0
10
0 1 2 0 0 8320 0 0 6 4 0 5
389 139
389 172
319 172
319 196
327 196
0 2 3 0 0 8192 0 0 7 3 0 5
400 205
400 159
321 159
321 148
329 148
3 1 3 0 0 4224 0 6 4 0 0 3
378 205
482 205
482 113
3 1 2 0 0 128 0 7 5 0 0 3
380 139
443 139
443 114
3 2 4 0 0 4224 0 8 6 0 0 4
255 209
319 209
319 214
327 214
3 1 5 0 0 4224 0 9 7 0 0 4
252 133
321 133
321 130
329 130
0 1 6 0 0 4224 0 0 2 8 0 4
193 170
117 170
117 169
108 169
1 2 6 0 0 0 0 8 9 0 0 4
204 200
193 200
193 142
201 142
1 2 7 0 0 8336 0 1 8 0 0 5
104 210
104 212
196 212
196 218
204 218
1 1 8 0 0 4224 0 3 9 0 0 4
109 123
193 123
193 124
201 124
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
464 42 501 66
474 50 490 66
2 QB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
429 43 458 67
439 51 447 67
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
51 194 80 218
61 202 69 218
1 R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
51 154 80 178
61 162 69 178
1 T
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
50 108 79 132
60 116 68 132
1 S
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
