CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 8 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
43032754 0
0
6 Title:
5 Name:
0
0
0
13
10 4-In NAND~
219 255 102 0 5 22
0 7 8 9 10 6
0
0 0 624 180
6 74LS20
-21 -40 21 -32
3 U5B
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
3277 0 0
2
42292.9 0
0
6 74LS48
188 597 413 0 14 29
0 21 22 23 24 32 33 20 19 18
17 16 15 14 34
0
0 0 4848 0
6 74LS48
-21 -76 21 -68
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4212 0 0
2
42292.9 5
0
9 Inverter~
13 269 480 0 2 22
0 11 10
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U7F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
4720 0 0
2
42292.9 2
0
9 Inverter~
13 293 478 0 2 22
0 12 9
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U7E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
5551 0 0
2
42292.9 1
0
6 74LS48
188 389 412 0 14 29
0 11 12 8 7 35 36 31 30 29
28 27 26 25 37
0
0 0 4848 0
6 74LS48
-21 -76 21 -68
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6986 0 0
2
42292.9 0
0
9 CC 7-Seg~
183 176 463 0 12 19
10 14 15 16 17 18 19 20 2 2
1 1 1
0
0 0 21088 0
7 AMBERCC
-77 -28 -28 -20
5 DISP1
-70 -15 -35 -7
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
8745 0 0
2
42292.8 2
0
9 CC 7-Seg~
183 71 464 0 16 19
10 25 26 27 28 29 30 31 2 2
1 1 0 1 1 0 1
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP2
34 -4 69 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
9592 0 0
2
42292.8 1
0
7 Ground~
168 169 588 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8748 0 0
2
42292.8 0
0
7 74LS161
96 141 129 0 14 29
0 5 4 3 38 39 40 41 5 6
42 11 12 8 7
0
0 0 4848 0
8 74LS161A
-24 -72 32 -64
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
7168 0 0
2
42292.8 0
0
7 74LS160
124 462 121 0 14 29
0 13 13 3 13 43 44 45 46 13
4 21 22 23 24
0
0 0 4848 0
8 74LS160A
-25 -61 31 -53
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
631 0 0
2
42292.8 0
0
7 Pulser~
4 300 37 0 10 12
0 47 48 3 49 0 0 5 5 2
8
0
0 0 4656 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9466 0 0
2
5.89727e-315 5.32571e-315
0
2 +V
167 81 23 0 1 3
0 5
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3266 0 0
2
5.89727e-315 5.46818e-315
0
2 +V
167 418 34 0 1 3
0 13
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7693 0 0
2
5.89727e-315 5.49538e-315
0
78
0 3 3 0 0 8320 0 0 9 70 0 5
385 112
385 269
47 269
47 111
109 111
2 10 4 0 0 12416 0 9 10 0 0 8
109 102
81 102
81 207
550 207
550 102
516 102
516 121
494 121
1 0 5 0 0 4096 0 12 0 0 13 2
81 32
81 55
9 5 6 0 0 4224 0 9 1 0 0 2
179 102
228 102
1 0 7 0 0 4096 0 1 0 0 9 2
279 115
312 115
2 1 8 0 0 4096 0 1 0 0 9 2
279 106
312 106
3 2 9 0 0 4096 0 1 0 0 9 2
279 97
312 97
4 3 10 0 0 4096 0 1 0 0 9 2
279 88
312 88
2 0 1 0 0 4128 0 0 0 0 0 2
312 72
312 128
11 3 11 0 0 4096 0 9 0 0 16 2
173 138
224 138
12 2 12 0 0 4096 0 9 0 0 16 2
173 147
224 147
13 1 8 0 0 4096 0 9 0 0 16 2
173 156
224 156
1 8 5 0 0 12416 0 9 9 0 0 6
109 93
81 93
81 55
191 55
191 93
179 93
0 9 13 0 0 4224 0 0 10 73 0 4
418 55
516 55
516 94
500 94
14 0 7 0 0 4096 0 9 0 0 16 2
173 165
224 165
1 0 1 0 0 32 0 0 0 0 0 2
224 122
224 171
13 0 14 0 0 4096 0 2 0 0 24 2
629 431
668 431
12 1 15 0 0 4096 0 2 0 0 24 2
629 422
668 422
11 2 16 0 0 4096 0 2 0 0 24 2
629 413
668 413
10 3 17 0 0 4096 0 2 0 0 24 2
629 404
668 404
9 4 18 0 0 4096 0 2 0 0 24 2
629 395
668 395
8 5 19 0 0 4096 0 2 0 0 24 2
629 386
668 386
7 6 20 0 0 4096 0 2 0 0 24 2
629 377
668 377
6 0 1 0 0 4256 0 0 0 0 0 2
668 369
668 440
3 1 21 0 0 4224 0 0 2 29 0 2
485 377
565 377
2 2 22 0 0 4224 0 0 2 29 0 2
485 386
565 386
1 3 23 0 0 4224 0 0 2 29 0 2
485 395
565 395
0 4 24 0 0 4224 0 0 2 29 0 2
485 404
565 404
4 0 1 0 0 32 0 0 0 0 0 2
485 360
485 409
2 3 10 0 0 4224 0 3 0 0 44 4
272 498
272 553
294 553
294 581
2 2 9 0 0 4224 0 4 0 0 44 4
296 496
296 542
303 542
303 581
0 1 11 0 0 4096 0 0 3 45 0 4
290 376
290 439
272 439
272 462
1 0 12 0 0 4096 0 4 0 0 46 2
296 460
296 385
13 0 25 0 0 4096 0 5 0 0 41 2
421 430
460 430
12 1 26 0 0 4096 0 5 0 0 41 2
421 421
460 421
11 2 27 0 0 4096 0 5 0 0 41 2
421 412
460 412
10 3 28 0 0 4096 0 5 0 0 41 2
421 403
460 403
9 4 29 0 0 4096 0 5 0 0 41 2
421 394
460 394
8 5 30 0 0 4096 0 5 0 0 41 2
421 385
460 385
7 6 31 0 0 4096 0 5 0 0 41 2
421 376
460 376
3 0 1 0 0 32 0 0 0 0 0 2
460 368
460 439
0 0 7 0 0 4224 0 0 0 48 44 2
323 403
323 581
1 0 8 0 0 4224 0 0 0 44 47 2
310 581
310 394
2 0 1 0 0 32 0 0 0 0 0 2
280 581
334 581
3 1 11 0 0 4224 0 0 5 49 0 2
275 376
357 376
2 2 12 0 0 4224 0 0 5 49 0 2
275 385
357 385
1 3 8 0 0 0 0 0 5 49 0 2
275 394
357 394
0 4 7 0 0 0 0 0 5 49 0 2
275 403
357 403
1 0 1 0 0 32 0 0 0 0 0 2
275 359
275 408
8 0 2 0 0 8192 0 7 0 0 53 3
92 500
92 519
112 519
8 0 2 0 0 8192 0 6 0 0 52 3
197 499
197 519
225 519
1 9 2 0 0 8320 0 8 6 0 0 4
169 582
225 582
225 421
176 421
9 1 2 0 0 0 0 7 8 0 0 4
71 422
112 422
112 582
169 582
1 0 14 0 0 4224 0 6 0 0 61 2
155 499
155 545
2 1 15 0 0 4224 0 6 0 0 61 2
161 499
161 545
3 2 16 0 0 4224 0 6 0 0 61 2
167 499
167 545
4 3 17 0 0 4224 0 6 0 0 61 2
173 499
173 545
5 4 18 0 0 4224 0 6 0 0 61 2
179 499
179 545
6 5 19 0 0 4224 0 6 0 0 61 2
185 499
185 545
7 6 20 0 0 4224 0 6 0 0 61 2
191 499
191 545
6 0 1 0 0 32 0 0 0 0 0 2
146 545
210 545
1 0 25 0 0 4224 0 7 0 0 69 2
50 500
50 546
2 1 26 0 0 4224 0 7 0 0 69 2
56 500
56 546
3 2 27 0 0 4224 0 7 0 0 69 2
62 500
62 546
4 3 28 0 0 4224 0 7 0 0 69 2
68 500
68 546
5 4 29 0 0 4224 0 7 0 0 69 2
74 500
74 546
6 5 30 0 0 4224 0 7 0 0 69 2
80 500
80 546
7 6 31 0 0 4224 0 7 0 0 69 2
86 500
86 546
3 0 1 0 0 32 0 0 0 0 0 2
41 546
105 546
3 3 3 0 0 128 0 11 10 0 0 4
324 28
385 28
385 112
430 112
1 0 13 0 0 0 0 10 0 0 73 2
430 94
418 94
2 0 13 0 0 0 0 10 0 0 73 2
430 103
418 103
1 4 13 0 0 128 0 13 10 0 0 3
418 43
418 121
424 121
11 3 21 0 0 0 0 10 0 0 78 2
494 130
538 130
12 2 22 0 0 0 0 10 0 0 78 2
494 139
538 139
13 1 23 0 0 0 0 10 0 0 78 2
494 148
538 148
14 0 24 0 0 0 0 10 0 0 78 2
494 157
538 157
4 0 1 0 0 32 0 0 0 0 0 2
538 116
538 165
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
