eNrtW+tzojoU/1cYvi7tABWKnbkfbGUtU18XH93OuuOwGFvm8nABb1/j/35PAHlYsHhdXW2zM81q
kpOT5PzyOL8TX+meYc1NzTccu+s6M+T6BvLoi1e6b1io7liaYeNvdflrbdDsj3tyv6+0Gz36wnfn
iKG7ziNya7ZmPnsGiE0100OLBUPLv+ZBm5D3/ZWeGXbfabjGhL6gWZqhvWfrp2N2Hc/AdSCTr7JP
PEsvfjD0lWPNHBvZvjc00COUqUgzQebWcMOOVSssx7M4lVj8feo61h19AXkM7Tv4kwSfcO43+gKq
4dzwE/RLlLDwOY/TfGE+ERalpTAIgLDEsbyENfMZzby0FOZTmqFyVjPHVlmxCklKtLqUrKa0xoJQ
GwQrwXgh5dn8LkN+LFyJx1uppISlUuNNCUtY+FzEYjCQMsJQORIGgXCyIuESZkomKxTGcyzmzLSY
N9OrNsZmEtnQWO8Kr2o+F8BCEve+maBiRjC07+pcVXNxlViYi4wEnauUG+2qhYO+SqX0ro411Chy
pfCc6BVT9g0X47vgWF0MQoAssRyyBDGrORQTyyFrda7D0UJ6xuWP+Yx7T1gqN2Ei9wYgYFGxHCxz
NOMxl1vHKWFYxyD94jgWVMH7hGJ7vmbr4Vaq8rC/vo5oua70a5dNeURfjGi8sY9oZkQ3lUu1pt6N
G2pn0A2Kgmx9uUGP/ecZCvI1OACc+6DUiNpva1ZYpvJRY1dyuyeP+3fdUA0bZMdf1eDrLD6Cgszv
r6PRiO5dd27HXbXTldX+Hc64wEnQzRGWgqSltMfDWnMgx8VsXHat1OtyOy4Ijqi4MNC/LFLlWjMu
6Q0urxT1aqD0x+1aK6kUV6gPWt1g0nJ7NGivCnYeLI+5CdIWTuOq2Y6DIZO+ZxpQk7515Sul1hwH
SrLi2Q5kyxj0hT3DiZhS0FeG8rhAT6v2rXBaU/Oj1INye26aieroxpCMK0+yoO91uXelKt2+0kns
piK4YQTQyp+GfCNlqqx2KanVVOqyqsp/DxRVrr+FyoJZA8QsoDZAYgYvewRiAfB48VQS8pHXR9Zs
W/CthVxGwe9E3Zag8+LLMeVDF5Gr+XMXUYZNTdC9ixB1hUzdmHsEkjuBZMFG2Ne53aIx1f4BgXFq
uJ5POe4EuRk06g6aTg3dgCOZ4HC/OOR3jEP+IDdFpDv2hADxwM5o27F2i8a0ggOCYxqBmk89Phj6
AzXTXHBAfOR61COCAvTku5ruo8kfAOaPwLVZsl1QDB7XE/wnVSunApQ8w2cee3kp3ypxn4Jrr+MG
bSjtXn/cu2tddppB4VdT8x4yNbz5zzrydNeYRbqgBeovCjsV1E3oddhBRdfxtbgKxwV5aasnPpmH
TIRnrpv1zcLCtEFwbgPZyDV0KtOpqWnMgtIv8C/UDrrt+5SPlzFAt6U9rTU5lMPFzKJ+ukj7h5ph
DpLSdNfxPMqNFJ+uwzk6AT8o8IbWIj7bxBqH5s2eEwM+s2UEZGnxlpDdpN7i0rplbpmb26Iz6pQX
3nd6IzBmCdgEkphKiwDJs4sFzdAdT2d3TxJgLaVoAqiYSxQUrTFRWq6wCpe/wKBFwzQdT3dmqHiR
vamVWT8sm7t+lp1dXSRvGlu/QNab7Jxfmuw8tFjDnuzBYlhLKYtBxY0sJkhSvCuesUK+0RquM4/a
zTVXqryMoZZ9fLObJc1sYyLMx0UDilaVyu2BeOMI8bYR8cYR4o0Qb4R4I8QbgSQh3gjxRog3QrwR
IBLi7eMRb+J5QrxxOybeuLXEW4E/Soi3z0a8JSwOF1EEja9zW98Dj4PVlCIKhpr+4amCIWMNmfmw
wNIFB8Bge3oALwtI1tMDg50cAuyWp8AM7wT/Oqav3Qf+Gf54aG7Z0eHw+oW5gb8W/DWuX4oIq3w4
Tn8fW4WT6lpMTg+Sspq66Ncc2fozBuQ1bFYvH+Va/McQuZmD1n3QPLTTS3FWwwHdig0bjnbNpGa4
gwlhRZiq/TIED8jXduuVZTQcEAAnmjWDOz41BbfLcQ/I7arwsdNV5U8LInuafjIMLxMnPWfu6mti
sj3DRkW+1wB8L4GCi5w9xV4YdYNP0fIO2PKuW+CCDZhprhNmTBCsfE2noiFQqSFsE0CsJGH5syiA
eLaHAOLZtgHEkuGkjxRE/IgRxE1chBIX8H0fgL8lvkTCi8caXixz/zkESG4SZSKRxeOLLB4LDjeK
MpHQ4vGFFo8FiP8zvkSCjMcaZDwsYBa5sefi/p7tU0f5ZH9NWG73McGtw5ZHFjmUuNUn+6qwB25A
II+LPz0vwJOXxcT1Jy+LCSSJ/09eFhP3n7wsJkAkTv+nflks7JMbaJHf85NnxWV/eRyTA5U9kAMV
Qg5sQg4I7Gd/NUDYAcIOEHaAQJKwA4QdIOwAYQcIEAk78PHYgcr+fncssBT50TFhB9azA8LKj44X
i/8ApHj3lw==