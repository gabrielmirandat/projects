* C:\Users\Marina\Desktop\exp5.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 20 14:54:14 2015



** Analysis setup **
.ac DEC 101 4.0K 400K


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "exp5.net"
.INC "exp5.als"


.probe


.END
