CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
43032754 0
0
6 Title:
5 Name:
0
0
0
48
13 Logic Switch~
5 44 502 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 NSCAR
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8838 0 0
2
42291 0
0
13 Logic Switch~
5 44 543 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
5 EWCAR
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7159 0 0
2
42291 1
0
9 2-In AND~
219 941 158 0 3 22
0 12 13 9
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
5812 0 0
2
42291 0
0
9 Inverter~
13 433 274 0 2 22
0 17 15
0
0 0 624 0
5 74F04
-50 -22 -15 -14
4 U16E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
331 0 0
2
42291 0
0
9 3-In AND~
219 529 274 0 4 22
0 16 15 18 14
0
0 0 624 0
6 74LS11
-23 21 19 29
3 U5A
-11 32 10 40
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 6 0
1 U
9604 0 0
2
42291 0
0
2 +V
167 415 38 0 1 3
0 19
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7518 0 0
2
42291 0
0
9 4-In NOR~
219 729 153 0 5 22
0 18 17 16 22 21
0
0 0 624 270
4 4002
30 3 58 11
4 U21A
30 -8 58 0
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 12 0
1 U
4832 0 0
2
42291 0
0
7 Ground~
168 414 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6798 0 0
2
42291 0
0
7 Ground~
168 96 189 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3336 0 0
2
42291 0
0
7 74LS160
124 462 121 0 14 29
0 19 19 21 23 2 2 2 2 19
67 58 59 12 13
0
0 0 4848 0
8 74LS160A
-25 -61 31 -53
2 U2
-8 -52 6 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
8370 0 0
2
42291 0
0
7 Ground~
168 140 366 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3910 0 0
2
42291 2
0
10 StopLight~
181 1122 503 0 12 13
0 7 6 3 0 0 0 0 0 0
0 0 1
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM2
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
316 0 0
2
42291 4
0
10 StopLight~
181 1120 401 0 10 13
0 8 5 4 0 0 0 0 0 0
1
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM1
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
536 0 0
2
42291 5
0
9 Inverter~
13 950 571 0 2 22
0 27 4
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U16D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
4460 0 0
2
42291 6
0
9 Inverter~
13 951 528 0 2 22
0 25 3
0
0 0 624 0
5 74F04
-50 -22 -15 -14
4 U16C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
3260 0 0
2
42291 7
0
10 2-In NAND~
219 956 446 0 3 22
0 29 24 5
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5156 0 0
2
42291 8
0
10 2-In NAND~
219 957 489 0 3 22
0 26 28 6
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3133 0 0
2
42291 9
0
2 +V
167 919 266 0 1 3
0 32
0
0 0 54256 0
3 10V
29 -11 50 -3
2 V8
13 -11 27 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5523 0 0
2
42291 10
0
10 8-In NAND~
219 957 392 0 9 19
0 32 32 32 31 30 29 24 27 7
0
0 0 624 0
6 74LS30
-21 -24 21 -16
3 U20
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
3746 0 0
2
42291 11
0
10 8-In NAND~
219 957 315 0 9 19
0 32 32 32 31 28 26 25 30 8
0
0 0 624 0
6 74LS30
-21 -24 21 -16
3 U19
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
5668 0 0
2
42291 12
0
7 Ground~
168 718 596 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5368 0 0
2
42291 13
0
2 +V
167 744 597 0 1 3
0 38
0
0 0 54256 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8293 0 0
2
42291 14
0
7 74LS138
19 790 535 0 14 29
0 35 34 33 38 2 2 31 28 26
25 30 29 24 27
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
3 U18
-11 -71 10 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3232 0 0
2
42291 15
0
7 Pulser~
4 67 411 0 10 12
0 68 69 11 70 0 0 5 5 2
7
0
0 0 4656 0
0
2 V2
-8 22 6 30
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6644 0 0
2
42291 16
0
2 +V
167 592 474 0 1 3
0 39
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4978 0 0
2
42291 17
0
7 Ground~
168 452 479 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9207 0 0
2
42291 18
0
9 Inverter~
13 602 505 0 2 22
0 37 36
0
0 0 624 180
5 74F04
13 -17 48 -9
4 U16B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
6998 0 0
2
42291 19
0
9 3-In AND~
219 640 559 0 4 22
0 35 34 33 37
0
0 0 624 0
6 74LS11
-23 21 19 29
4 U15C
-14 32 14 40
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 10 0
1 U
3175 0 0
2
42291 20
0
7 74LS161
96 542 532 0 14 29
0 40 40 11 71 72 73 74 39 36
75 76 35 34 33
0
0 0 4848 0
8 74LS161A
-27 -71 29 -63
3 U17
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3378 0 0
2
42291 21
0
8 2-In OR~
219 285 534 0 3 22
0 9 42 48
0
0 0 624 0
6 74LS32
5 -30 47 -22
4 U14B
-26 -29 2 -21
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
922 0 0
2
42291 22
0
8 2-In OR~
219 285 570 0 3 22
0 9 41 47
0
0 0 624 0
6 74LS32
5 19 47 27
4 U14A
-23 20 5 28
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
6891 0 0
2
42291 23
0
2 +V
167 343 602 0 1 3
0 49
0
0 0 54256 180
3 10V
9 -3 30 5
2 V5
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5407 0 0
2
42291 24
0
7 74LS151
20 399 534 0 14 29
0 49 49 49 48 49 49 49 47 2
35 34 33 40 77
0
0 0 4848 0
7 74LS151
-24 -72 25 -64
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7349 0 0
2
42291 25
0
9 3-In AND~
219 212 579 0 4 22
0 46 45 10 41
0
0 0 624 0
6 74LS11
-47 17 -5 25
4 U15B
2 17 30 25
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 10 0
1 U
3919 0 0
2
42291 27
0
9 3-In AND~
219 212 543 0 4 22
0 43 44 10 42
0
0 0 624 0
6 74LS11
-40 -26 2 -18
4 U15A
3 -26 31 -18
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 10 0
1 U
9747 0 0
2
42291 28
0
9 Inverter~
13 95 522 0 2 22
0 45 43
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
5310 0 0
2
42291 29
0
9 Inverter~
13 96 471 0 2 22
0 44 46
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
4318 0 0
2
42291 30
0
2 +V
167 102 45 0 1 3
0 20
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3917 0 0
2
42291 31
0
6 74LS48
188 1022 79 0 14 29
0 58 59 12 13 78 79 57 56 55
54 53 52 51 80
0
0 0 4848 0
6 74LS48
-21 -76 21 -68
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7930 0 0
2
42291 41
0
6 74LS48
188 814 78 0 14 29
0 22 16 17 18 81 82 66 65 64
63 62 61 60 83
0
0 0 4848 0
6 74LS48
-21 -76 21 -68
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6128 0 0
2
42291 46
0
9 CC 7-Seg~
183 88 244 0 15 19
10 51 52 53 54 55 56 57 2 2
1 1 1 1 1 1
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP2
34 -4 69 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
7346 0 0
2
42291 48
0
9 CC 7-Seg~
183 193 243 0 12 19
10 60 61 62 63 64 65 66 2 2
0 1 1
0
0 0 21088 0
7 AMBERCC
-77 -28 -28 -20
5 DISP1
-70 -15 -35 -7
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
8577 0 0
2
42291 49
0
7 74LS160
124 145 139 0 14 29
0 20 20 11 23 2 2 2 2 20
84 22 16 17 18
0
0 0 4848 0
8 74LS160A
-25 -61 31 -53
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3372 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 793 232 0 1 2
10 9
0
0 0 53856 0
6 100MEG
11 -9 53 -1
6 TMLONG
-10 -21 32 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3741 0 0
2
5.89727e-315 5.30499e-315
0
2 +V
167 612 200 0 1 3
0 50
0
0 0 54256 0
3 10V
8 -2 29 6
2 V4
12 8 26 16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5813 0 0
2
5.89727e-315 5.32571e-315
0
14 Logic Display~
6 749 232 0 1 2
10 10
0
0 0 53856 0
6 100MEG
-51 -7 -9 1
7 TMSHORT
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3213 0 0
2
5.89727e-315 5.34643e-315
0
10 2-In NAND~
219 264 38 0 3 22
0 8 7 23
0
0 0 624 0
4 7400
-15 -36 13 -28
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3694 0 0
2
5.89727e-315 5.3568e-315
0
5 7474~
219 612 292 0 6 22
0 50 50 14 23 85 10
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
4327 0 0
2
42291 50
0
164
3 0 11 0 0 8192 0 43 0 0 82 5
113 130
34 130
34 369
109 369
109 402
3 1 9 0 0 8192 0 3 44 0 0 6
939 181
939 206
865 206
865 276
793 276
793 250
1 0 12 0 0 4096 0 3 0 0 123 2
948 136
948 61
2 0 13 0 0 4096 0 3 0 0 124 2
930 136
930 70
4 3 14 0 0 4224 0 5 48 0 0 2
550 274
588 274
2 2 15 0 0 4224 0 4 5 0 0 2
454 274
505 274
1 2 16 0 0 8320 0 5 0 0 10 3
505 265
505 261
341 261
1 1 17 0 0 12288 0 0 4 10 0 4
341 276
356 276
356 274
418 274
3 0 18 0 0 8336 0 5 0 0 10 3
505 283
505 292
341 292
1 0 1 0 0 4128 0 0 0 0 0 2
341 250
341 299
9 0 19 0 0 12416 0 10 0 0 13 4
500 94
514 94
514 55
415 55
0 2 19 0 0 0 0 0 10 13 0 3
415 94
415 103
430 103
1 1 19 0 0 0 0 6 10 0 0 3
415 47
415 94
430 94
0 9 20 0 0 4224 0 0 43 16 0 4
102 70
199 70
199 112
183 112
0 2 20 0 0 0 0 0 43 16 0 3
102 111
102 121
113 121
1 1 20 0 0 0 0 38 43 0 0 3
102 54
102 112
113 112
3 5 21 0 0 12416 0 10 7 0 0 7
430 112
388 112
388 184
710 184
710 195
735 195
735 186
1 0 18 0 0 0 0 7 0 0 137 2
748 130
748 69
2 0 17 0 0 4096 0 7 0 0 136 2
739 130
739 60
3 0 16 0 0 0 0 7 0 0 135 2
730 130
730 51
4 0 22 0 0 4224 0 7 0 0 134 2
721 130
721 42
0 5 2 0 0 8192 0 0 10 23 0 3
414 139
414 130
430 130
0 6 2 0 0 0 0 0 10 24 0 3
414 149
414 139
430 139
0 7 2 0 0 0 0 0 10 25 0 3
414 157
414 148
430 148
1 8 2 0 0 0 0 8 10 0 0 3
414 165
414 157
430 157
0 5 2 0 0 8192 0 0 43 27 0 3
96 157
96 148
113 148
0 6 2 0 0 0 0 0 43 28 0 3
96 167
96 157
113 157
0 7 2 0 0 0 0 0 43 29 0 3
96 175
96 166
113 166
1 8 2 0 0 0 0 9 43 0 0 3
96 183
96 175
113 175
0 4 23 0 0 16512 0 0 48 31 0 6
401 120
401 193
281 193
281 386
612 386
612 304
0 4 23 0 0 0 0 0 10 32 0 4
303 62
401 62
401 121
424 121
3 4 23 0 0 0 0 47 43 0 0 6
291 38
303 38
303 62
91 62
91 139
107 139
2 0 24 0 0 4096 0 16 0 0 56 2
932 455
887 455
8 0 2 0 0 8192 0 41 0 0 37 3
109 280
109 299
129 299
8 0 2 0 0 8192 0 42 0 0 36 3
214 279
214 299
242 299
1 9 2 0 0 8320 0 11 42 0 0 4
140 360
242 360
242 201
193 201
9 1 2 0 0 0 0 41 11 0 0 4
88 202
129 202
129 360
140 360
3 2 6 0 0 12416 0 17 12 0 0 4
984 489
1025 489
1025 503
1106 503
0 1 7 0 0 8320 0 0 12 44 0 4
991 392
1074 392
1074 489
1106 489
0 1 8 0 0 4224 0 0 13 45 0 4
994 315
1084 315
1084 387
1104 387
2 1 7 0 0 0 0 47 0 0 43 2
240 47
164 47
1 0 8 0 0 0 0 47 0 0 43 2
240 29
164 29
7 0 1 0 0 32 0 0 0 0 0 2
164 20
164 55
9 1 7 0 0 0 0 19 0 0 46 4
984 392
991 392
991 349
1025 349
9 0 8 0 0 0 0 20 0 0 46 4
984 315
994 315
994 335
1025 335
7 0 1 0 0 32 0 0 0 0 0 2
1025 322
1025 361
1 0 25 0 0 4096 0 15 0 0 67 2
936 528
863 528
1 0 26 0 0 4096 0 17 0 0 68 2
933 480
854 480
1 0 27 0 0 4096 0 14 0 0 55 2
935 571
894 571
2 0 28 0 0 4096 0 17 0 0 69 2
933 498
845 498
1 0 29 0 0 4096 0 16 0 0 57 2
932 437
879 437
2 3 4 0 0 16512 0 14 13 0 0 6
971 571
1062 571
1062 561
1087 561
1087 415
1104 415
2 3 3 0 0 4224 0 15 12 0 0 4
972 528
1062 528
1062 517
1106 517
3 2 5 0 0 4224 0 16 13 0 0 4
983 446
1059 446
1059 401
1104 401
14 8 27 0 0 8320 0 23 19 0 0 4
828 571
896 571
896 424
933 424
13 7 24 0 0 8320 0 23 19 0 0 4
828 562
887 562
887 415
933 415
12 6 29 0 0 8320 0 23 19 0 0 4
828 553
879 553
879 406
933 406
5 0 30 0 0 4096 0 19 0 0 66 2
933 397
871 397
4 0 31 0 0 4096 0 19 0 0 70 2
933 388
837 388
0 3 32 0 0 4096 0 0 19 61 0 2
919 379
933 379
0 2 32 0 0 0 0 0 19 62 0 5
919 370
919 379
919 379
919 370
933 370
0 1 32 0 0 4224 0 0 19 63 0 5
919 301
919 370
919 370
919 361
933 361
0 3 32 0 0 0 0 0 20 64 0 3
919 293
919 302
933 302
0 2 32 0 0 0 0 0 20 65 0 3
919 283
919 293
933 293
1 1 32 0 0 0 0 18 20 0 0 3
919 275
919 284
933 284
11 8 30 0 0 8320 0 23 20 0 0 4
828 544
871 544
871 347
933 347
10 7 25 0 0 8320 0 23 20 0 0 4
828 535
863 535
863 338
933 338
9 6 26 0 0 8320 0 23 20 0 0 4
828 526
854 526
854 329
933 329
8 5 28 0 0 8320 0 23 20 0 0 4
828 517
845 517
845 320
933 320
7 4 31 0 0 8320 0 23 20 0 0 4
828 508
837 508
837 311
933 311
0 12 33 0 0 8320 0 0 33 76 0 5
608 568
608 601
452 601
452 534
431 534
0 11 34 0 0 8320 0 0 33 75 0 5
601 559
601 593
461 593
461 525
431 525
0 10 35 0 0 8192 0 0 33 74 0 5
594 550
594 585
470 585
470 516
431 516
0 1 35 0 0 8320 0 0 23 88 0 5
594 550
594 522
719 522
719 508
758 508
0 2 34 0 0 0 0 0 23 89 0 5
601 559
601 530
727 530
727 517
758 517
0 3 33 0 0 0 0 0 23 87 0 5
608 568
608 539
735 539
735 526
758 526
2 9 36 0 0 12416 0 27 29 0 0 4
587 505
588 505
588 505
580 505
1 4 37 0 0 8320 0 27 28 0 0 4
623 505
673 505
673 559
661 559
0 5 2 0 0 0 0 0 23 80 0 3
718 572
718 562
752 562
1 6 2 0 0 0 0 21 23 0 0 3
718 590
718 571
752 571
1 4 38 0 0 4224 0 22 23 0 0 3
744 582
744 553
758 553
3 3 11 0 0 12416 0 29 24 0 0 4
510 514
494 514
494 402
91 402
8 1 39 0 0 8320 0 29 25 0 0 3
580 496
592 496
592 483
2 0 40 0 0 4096 0 29 0 0 85 2
510 505
475 505
13 1 40 0 0 8320 0 33 29 0 0 4
431 561
475 561
475 496
510 496
9 1 2 0 0 0 0 33 26 0 0 3
437 507
452 507
452 487
3 14 33 0 0 0 0 28 29 0 0 2
616 568
574 568
12 1 35 0 0 0 0 29 28 0 0 2
574 550
616 550
13 2 34 0 0 0 0 29 28 0 0 2
574 559
616 559
4 2 41 0 0 4224 0 34 31 0 0 2
233 579
272 579
4 2 42 0 0 4224 0 35 30 0 0 2
233 543
272 543
2 1 43 0 0 12416 0 36 35 0 0 4
116 522
138 522
138 534
188 534
0 2 44 0 0 4224 0 0 35 109 0 4
66 489
164 489
164 543
188 543
0 3 10 0 0 4096 0 0 34 95 0 3
173 552
173 588
188 588
0 3 10 0 0 8320 0 0 35 110 0 5
749 320
749 444
173 444
173 552
188 552
0 2 45 0 0 8320 0 0 34 108 0 3
66 543
66 579
188 579
2 1 46 0 0 8320 0 37 34 0 0 4
117 471
156 471
156 570
188 570
0 1 9 0 0 0 0 0 31 99 0 3
263 523
263 561
272 561
0 1 9 0 0 8320 0 0 30 2 0 5
793 276
793 414
263 414
263 525
272 525
3 8 47 0 0 4224 0 31 33 0 0 2
318 570
367 570
3 4 48 0 0 4224 0 30 33 0 0 2
318 534
367 534
3 0 49 0 0 4096 0 33 0 0 104 2
367 525
343 525
2 0 49 0 0 0 0 33 0 0 104 2
367 516
343 516
0 1 49 0 0 4224 0 0 33 105 0 3
343 543
343 507
367 507
0 5 49 0 0 0 0 0 33 106 0 3
343 553
343 543
367 543
0 6 49 0 0 0 0 0 33 107 0 3
343 561
343 552
367 552
1 7 49 0 0 0 0 32 33 0 0 3
343 587
343 561
367 561
1 1 45 0 0 0 0 2 36 0 0 4
56 543
67 543
67 522
80 522
1 1 44 0 0 0 0 1 37 0 0 4
56 502
66 502
66 471
81 471
6 1 10 0 0 0 0 48 46 0 0 5
636 256
675 256
675 320
749 320
749 250
2 0 50 0 0 12416 0 48 0 0 112 4
588 256
575 256
575 220
612 220
1 1 50 0 0 0 0 45 48 0 0 2
612 209
612 229
13 0 51 0 0 4096 0 39 0 0 120 2
1054 97
1093 97
12 1 52 0 0 4096 0 39 0 0 120 2
1054 88
1093 88
11 2 53 0 0 4096 0 39 0 0 120 2
1054 79
1093 79
10 3 54 0 0 4096 0 39 0 0 120 2
1054 70
1093 70
9 4 55 0 0 4096 0 39 0 0 120 2
1054 61
1093 61
8 5 56 0 0 4096 0 39 0 0 120 2
1054 52
1093 52
7 6 57 0 0 4096 0 39 0 0 120 2
1054 43
1093 43
6 0 1 0 0 4256 0 0 0 0 0 2
1093 35
1093 106
3 1 58 0 0 4224 0 0 39 125 0 2
910 43
990 43
2 2 59 0 0 4224 0 0 39 125 0 2
910 52
990 52
1 3 12 0 0 4224 0 0 39 125 0 2
910 61
990 61
0 4 13 0 0 4224 0 0 39 125 0 2
910 70
990 70
4 0 1 0 0 32 0 0 0 0 0 2
910 26
910 75
13 0 60 0 0 4096 0 40 0 0 133 2
846 96
885 96
12 1 61 0 0 4096 0 40 0 0 133 2
846 87
885 87
11 2 62 0 0 4096 0 40 0 0 133 2
846 78
885 78
10 3 63 0 0 4096 0 40 0 0 133 2
846 69
885 69
9 4 64 0 0 4096 0 40 0 0 133 2
846 60
885 60
8 5 65 0 0 4096 0 40 0 0 133 2
846 51
885 51
7 6 66 0 0 4096 0 40 0 0 133 2
846 42
885 42
3 0 1 0 0 32 0 0 0 0 0 2
885 34
885 105
3 1 22 0 0 128 0 0 40 138 0 2
700 42
782 42
2 2 16 0 0 128 0 0 40 138 0 2
700 51
782 51
1 3 17 0 0 4224 0 0 40 138 0 2
700 60
782 60
0 4 18 0 0 0 0 0 40 138 0 2
700 69
782 69
1 0 1 0 0 32 0 0 0 0 0 2
700 25
700 74
1 0 60 0 0 4224 0 42 0 0 146 2
172 279
172 325
2 1 61 0 0 4224 0 42 0 0 146 2
178 279
178 325
3 2 62 0 0 4224 0 42 0 0 146 2
184 279
184 325
4 3 63 0 0 4224 0 42 0 0 146 2
190 279
190 325
5 4 64 0 0 4224 0 42 0 0 146 2
196 279
196 325
6 5 65 0 0 4224 0 42 0 0 146 2
202 279
202 325
7 6 66 0 0 4224 0 42 0 0 146 2
208 279
208 325
3 0 1 0 0 32 0 0 0 0 0 2
163 325
227 325
1 0 51 0 0 4224 0 41 0 0 154 2
67 280
67 326
2 1 52 0 0 4224 0 41 0 0 154 2
73 280
73 326
3 2 53 0 0 4224 0 41 0 0 154 2
79 280
79 326
4 3 54 0 0 4224 0 41 0 0 154 2
85 280
85 326
5 4 55 0 0 4224 0 41 0 0 154 2
91 280
91 326
6 5 56 0 0 4224 0 41 0 0 154 2
97 280
97 326
7 6 57 0 0 4224 0 41 0 0 154 2
103 280
103 326
6 0 1 0 0 32 0 0 0 0 0 2
58 326
122 326
11 3 58 0 0 0 0 10 0 0 159 2
494 130
538 130
12 2 59 0 0 0 0 10 0 0 159 2
494 139
538 139
13 1 12 0 0 0 0 10 0 0 159 2
494 148
538 148
14 0 13 0 0 0 0 10 0 0 159 2
494 157
538 157
4 0 1 0 0 32 0 0 0 0 0 2
538 116
538 165
11 3 22 0 0 0 0 43 0 0 164 2
177 148
220 148
12 2 16 0 0 0 0 43 0 0 164 2
177 157
220 157
13 1 17 0 0 0 0 43 0 0 164 2
177 166
220 166
14 0 18 0 0 0 0 43 0 0 164 2
177 175
220 175
1 0 1 0 0 32 0 0 0 0 0 2
220 134
220 183
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
988 512 1047 528
988 512 1047 528
7 EWGREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
989 555 1048 571
989 555 1048 571
7 NSGREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 8
986 430 1053 446
986 430 1053 446
8 NSYELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 8
991 473 1058 489
991 473 1058 489
8 EWYELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
1001 376 1044 392
1001 376 1044 392
5 EWRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
992 299 1035 315
992 299 1035 315
5 NSRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
185 31 228 47
185 31 228 47
5 EWRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
188 13 231 29
188 13 231 29
5 NSRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 6
678 398 729 414
678 398 729 414
6 TMLONG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
676 304 735 320
676 304 735 320
7 TMSHORT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
