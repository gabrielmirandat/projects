CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
84 216 630 550
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 C:\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
252 312 365 409
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 58 80 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8495 0 0
2
42183 0
0
13 Logic Switch~
5 196 47 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
398 0 0
2
42183 0
0
13 Logic Switch~
5 195 225 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3192 0 0
2
42183 0
0
13 Logic Switch~
5 60 125 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3665 0 0
2
42183 0
0
13 Logic Switch~
5 64 179 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6514 0 0
2
42183 0
0
14 Logic Display~
6 378 67 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3703 0 0
2
42183 0
0
14 Logic Display~
6 346 69 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8955 0 0
2
42183 0
0
10 3-In NAND~
219 259 167 0 4 22
0 2 4 7 3
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 2 0
1 U
4449 0 0
2
42183 0
0
10 3-In NAND~
219 258 95 0 4 22
0 6 5 3 2
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
3268 0 0
2
42183 0
0
10 2-In NAND~
219 137 171 0 3 22
0 8 9 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5679 0 0
2
42183 0
0
10 2-In NAND~
219 137 93 0 3 22
0 10 8 5
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3376 0 0
2
42183 0
0
12
0 1 2 0 0 8192 0 0 8 4 0 5
285 95
285 131
227 131
227 158
235 158
0 3 3 0 0 8192 0 0 9 3 0 5
296 167
296 115
226 115
226 104
234 104
4 1 3 0 0 4224 0 8 6 0 0 3
286 167
378 167
378 85
4 1 2 0 0 4224 0 9 7 0 0 3
285 95
346 95
346 87
3 2 4 0 0 4224 0 10 8 0 0 4
164 171
227 171
227 167
235 167
3 2 5 0 0 4224 0 11 9 0 0 4
164 93
226 93
226 95
234 95
1 1 6 0 0 8320 0 2 9 0 0 4
208 47
226 47
226 86
234 86
1 3 7 0 0 8320 0 3 8 0 0 4
207 225
227 225
227 176
235 176
0 1 8 0 0 4096 0 0 4 10 0 2
105 125
72 125
1 2 8 0 0 8320 0 10 11 0 0 4
113 162
105 162
105 102
113 102
1 2 9 0 0 4224 0 5 10 0 0 4
76 179
105 179
105 180
113 180
1 1 10 0 0 8320 0 1 11 0 0 5
70 80
70 79
105 79
105 84
113 84
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
129 227 238 251
139 235 227 251
11 Clear barra
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
93 -2 210 22
103 6 199 22
12 Preset barra
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
359 22 396 46
369 30 385 46
2 QB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
329 20 358 44
339 28 347 44
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
26 115 55 139
36 123 44 139
1 T
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
31 167 60 191
41 175 49 191
1 R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
23 61 52 85
33 69 41 85
1 S
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
