CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
23 C:\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9469970 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 53 116 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5779 0 0
2
42181.9 0
0
13 Logic Switch~
5 34 229 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9443 0 0
2
42181.9 1
0
9 2-In NOR~
219 250 216 0 3 22
0 4 2 5
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8374 0 0
2
5.89713e-315 5.30499e-315
0
9 2-In NOR~
219 254 131 0 3 22
0 3 5 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4469 0 0
2
5.89713e-315 5.32571e-315
0
14 Logic Display~
6 393 104 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7424 0 0
2
42181.9 2
0
14 Logic Display~
6 350 106 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7305 0 0
2
42181.9 3
0
7
0 2 2 0 0 8320 0 0 3 3 0 3
116 234
116 225
237 225
1 1 3 0 0 4224 0 1 4 0 0 4
65 116
180 116
180 122
241 122
1 0 2 0 0 0 0 2 0 0 0 4
46 229
57 229
57 234
123 234
1 0 4 0 0 12416 0 3 0 0 7 5
237 207
219 207
219 179
304 179
304 134
2 0 5 0 0 12416 0 4 0 0 6 5
241 140
218 140
218 165
313 165
313 212
3 1 5 0 0 0 0 3 5 0 0 5
289 216
313 216
313 212
393 212
393 122
3 1 4 0 0 0 0 4 6 0 0 5
293 131
304 131
304 134
350 134
350 124
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
-1 213 28 237
9 221 17 237
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
10 92 39 116
20 100 28 116
1 R
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
376 55 413 79
386 63 402 79
2 QB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
335 58 364 82
345 66 353 82
1 Q
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
