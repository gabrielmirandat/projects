CircuitMaker Text
5.6
Probes: 1
rd2[i]
Transient Analysis
0 560 388 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
259 95 1274 632
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
427 191 540 288
1083744434 0
0
6 Title:
5 Name:
0
0
0
23
9 V Source~
197 283 436 0 2 5
0 5 2
0
0 0 17248 0
3 10V
13 0 34 8
3 Vs3
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
6369 0 0
2
42275.8 0
0
7 Ground~
168 366 528 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
42275.8 1
0
9 V Source~
197 475 206 0 2 5
0 9 2
0
0 0 17248 0
3 10V
13 0 34 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
7100 0 0
2
42275.8 2
0
7 Ground~
168 558 306 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
42275.8 3
0
7 Ground~
168 162 296 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
42275.8 4
0
9 V Source~
197 79 204 0 2 5
0 13 2
0
0 0 17248 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
961 0 0
2
42275.8 5
0
9 Resistor~
219 473 407 0 2 5
0 4 5
0
0 0 864 90
2 1k
8 0 22 8
3 Rb2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
42275.8 6
0
9 Resistor~
219 560 406 0 2 5
0 3 5
0
0 0 864 90
4 4700
3 0 31 8
3 Rd2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
42275.8 7
0
9 Resistor~
219 521 452 0 2 5
0 3 4
0
0 0 864 180
3 100
-10 -14 11 -6
3 Rf2
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
42275.8 8
0
9 Resistor~
219 474 491 0 3 5
0 2 4 -1
0
0 0 864 90
4 4700
1 0 29 8
3 Re2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
42275.8 9
0
9 Resistor~
219 560 493 0 3 5
0 2 3 -1
0
0 0 864 90
2 1k
8 0 22 8
3 Rc2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
42275.8 10
0
9 Resistor~
219 549 138 0 2 5
0 9 7
0
0 0 864 0
4 2011
-14 -14 14 -6
3 Ra1
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
42275.8 11
0
9 Resistor~
219 665 177 0 2 5
0 8 7
0
0 0 864 90
4 1035
1 0 29 8
3 Rb1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
42275.8 12
0
9 Resistor~
219 754 262 0 3 5
0 2 6 -1
0
0 0 864 90
4 4700
3 0 31 8
3 Rd1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9424 0 0
2
42275.8 13
0
9 Resistor~
219 713 222 0 2 5
0 6 8
0
0 0 864 180
3 100
-10 -14 11 -6
3 Rf1
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
42275.8 14
0
9 Resistor~
219 666 261 0 3 5
0 2 8 -1
0
0 0 864 90
4 4700
1 0 29 8
3 Re1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
42275.8 15
0
9 Resistor~
219 754 172 0 2 5
0 6 7
0
0 0 864 90
4 1035
1 0 29 8
3 Rc1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
42275.8 16
0
9 Resistor~
219 356 261 0 3 5
0 2 10 -1
0
0 0 864 90
4 1035
1 0 29 8
2 Rc
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66269076
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
42275.8 17
0
9 Resistor~
219 270 259 0 3 5
0 2 11 -1
0
0 0 864 90
4 4700
1 0 29 8
2 Re
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66269956
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
42275.8 18
0
9 Resistor~
219 317 220 0 2 5
0 10 11
0
0 0 864 180
3 100
-10 -14 11 -6
2 Rf
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 70
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
42275.8 19
0
9 Resistor~
219 356 174 0 2 5
0 10 12
0
0 0 864 90
4 4700
3 0 31 8
2 Rd
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 38
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
42275.8 20
0
9 Resistor~
219 269 175 0 2 5
0 11 12
0
0 0 864 90
4 1035
1 0 29 8
2 Rb
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
5283 0 0
2
42275.8 21
0
9 Resistor~
219 153 136 0 2 5
0 13 12
0
0 0 864 0
4 2011
-14 -14 14 -6
2 Ra
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 70
82 0 0 0 1 0 0 0
1 R
6874 0 0
2
42275.8 22
0
29
1 0 2 0 0 4096 0 10 0 0 2 2
474 509
474 522
1 1 2 0 0 4224 0 2 11 0 0 3
366 522
560 522
560 511
2 1 2 0 0 0 0 1 2 0 0 3
283 457
283 522
366 522
1 0 3 0 0 4096 0 9 0 0 5 2
539 452
560 452
1 2 3 0 0 4224 0 8 11 0 0 2
560 424
560 475
2 0 4 0 0 4096 0 9 0 0 7 2
503 452
474 452
1 2 4 0 0 8320 0 7 10 0 0 3
473 425
474 425
474 473
2 0 5 0 0 4096 0 7 0 0 9 2
473 389
473 368
1 2 5 0 0 8320 0 1 8 0 0 4
283 415
283 368
560 368
560 388
0 1 2 0 0 0 0 0 14 13 0 3
666 300
754 300
754 280
0 2 6 0 0 8192 0 0 14 15 0 3
753 222
754 222
754 244
0 2 7 0 0 4096 0 0 17 18 0 3
665 138
754 138
754 154
1 1 2 0 0 0 0 16 4 0 0 3
666 279
666 300
558 300
2 1 2 0 0 0 0 3 4 0 0 3
475 227
475 300
558 300
1 1 6 0 0 8320 0 15 17 0 0 3
731 222
754 222
754 190
2 0 8 0 0 4096 0 15 0 0 17 2
695 222
666 222
1 2 8 0 0 8320 0 13 16 0 0 3
665 195
666 195
666 243
2 2 7 0 0 8320 0 13 12 0 0 3
665 159
665 138
567 138
1 1 9 0 0 8320 0 3 12 0 0 3
475 185
475 138
531 138
1 0 2 0 0 0 0 19 0 0 21 2
270 277
270 290
1 1 2 0 0 0 0 5 18 0 0 3
162 290
356 290
356 279
2 1 2 0 0 0 0 6 5 0 0 3
79 225
79 290
162 290
1 0 10 0 0 4096 0 20 0 0 24 2
335 220
356 220
1 2 10 0 0 4224 0 21 18 0 0 2
356 192
356 243
2 0 11 0 0 4096 0 20 0 0 26 2
299 220
270 220
1 2 11 0 0 8320 0 22 19 0 0 3
269 193
270 193
270 241
2 0 12 0 0 4096 0 22 0 0 28 2
269 157
269 136
2 2 12 0 0 4224 0 23 21 0 0 3
171 136
356 136
356 156
1 1 13 0 0 8320 0 6 23 0 0 3
79 183
79 136
135 136
0
0
17 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
