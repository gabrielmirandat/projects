CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 284 114 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
42180.5 0
0
13 Logic Switch~
5 283 232 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
2 Ai
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
42180.5 0
0
13 Logic Switch~
5 284 171 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 Bi
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
42180.5 0
0
14 Logic Display~
6 693 185 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Si
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
42180.5 0
0
14 Logic Display~
6 673 137 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
4 Cout
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
42180.5 0
0
9 Inverter~
13 423 203 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
5572 0 0
2
42180.5 0
0
7 Ground~
168 403 356 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8901 0 0
2
42180.5 0
0
2 +V
167 405 33 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
42180.5 0
0
7 74LS153
119 508 171 0 14 29
0 8 7 7 2 9 3 7 6 6
7 2 2 5 4
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 0 0 0 0
1 U
4747 0 0
2
42180.5 0
0
15
1 6 3 0 0 12416 0 2 9 0 0 4
295 232
325 232
325 180
476 180
14 1 4 0 0 4224 0 9 4 0 0 3
540 198
693 198
693 203
13 1 5 0 0 4224 0 9 5 0 0 5
540 153
672 153
672 149
673 149
673 155
12 0 2 0 0 4096 0 9 0 0 5 2
546 216
579 216
11 0 2 0 0 8192 0 9 0 0 9 4
546 135
579 135
579 277
461 277
0 9 6 0 0 8320 0 0 9 7 0 3
452 203
452 207
476 207
2 8 6 0 0 0 0 6 9 0 0 4
444 203
453 203
453 198
476 198
0 1 7 0 0 8192 0 0 6 14 0 3
402 204
402 203
408 203
1 4 2 0 0 12416 0 7 9 0 0 5
403 350
403 317
461 317
461 162
476 162
1 1 8 0 0 8320 0 8 9 0 0 4
405 42
461 42
461 135
476 135
2 0 7 0 0 4096 0 9 0 0 14 2
476 144
402 144
3 0 7 0 0 0 0 9 0 0 14 2
476 153
402 153
7 0 7 0 0 0 0 9 0 0 14 2
476 189
402 189
1 10 7 0 0 8320 0 1 9 0 0 4
296 114
402 114
402 216
476 216
1 5 9 0 0 4224 0 3 9 0 0 2
296 171
476 171
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
