CircuitMaker Text
5.6
Probes: 1
C1_2
Transient Analysis
0 437 87 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
35
9 Inductor~
219 639 525 0 2 5
0 21 22
0
0 0 832 0
6 1.05mH
-21 -17 21 -9
2 L5
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
5130 0 0
2
42325.4 0
0
9 Inductor~
219 638 391 0 2 5
0 21 22
0
0 0 832 0
6 1.05mH
-21 -17 21 -9
2 L6
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
391 0 0
2
42325.4 0
0
9 Inductor~
219 628 240 0 2 5
0 21 22
0
0 0 832 0
6 1.05mH
-21 -17 21 -9
2 L7
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3124 0 0
2
42325.4 0
0
9 Inductor~
219 310 523 0 2 5
0 21 22
0
0 0 832 0
6 1.05mH
-21 -17 21 -9
2 L4
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3421 0 0
2
42325.4 0
0
9 Inductor~
219 310 391 0 2 5
0 21 22
0
0 0 832 0
6 1.05mH
-21 -17 21 -9
2 L3
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
8157 0 0
2
42325.4 0
0
10 Capacitor~
219 676 563 0 2 5
0 2 22
0
0 0 832 90
8 0.9272nF
-6 0 50 8
2 C5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5572 0 0
2
42325.4 0
0
10 Capacitor~
219 676 429 0 2 5
0 2 22
0
0 0 832 90
8 0.9272nF
-6 0 50 8
2 C6
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8901 0 0
2
42325.4 0
0
10 Capacitor~
219 667 277 0 2 5
0 2 22
0
0 0 832 90
8 0.9272nF
-6 0 50 8
2 C7
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7361 0 0
2
42325.4 0
0
10 Capacitor~
219 350 563 0 2 5
0 2 22
0
0 0 832 90
8 0.9272nF
-6 0 50 8
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4747 0 0
2
42325.4 0
0
10 Capacitor~
219 349 430 0 2 5
0 2 22
0
0 0 832 90
8 0.9272nF
-6 0 50 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
972 0 0
2
42325.4 0
0
10 Capacitor~
219 341 277 0 2 5
0 2 22
0
0 0 832 90
8 0.9272nF
-6 0 50 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3472 0 0
2
42325.4 0
0
11 Signal Gen~
195 497 422 0 64 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V6
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.89731e-315 5.4086e-315
0
7 Ground~
168 608 482 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.89731e-315 5.40342e-315
0
7 Ground~
168 608 616 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.89731e-315 5.39824e-315
0
11 Signal Gen~
195 497 556 0 64 64
0 5 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V5
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
5.89731e-315 5.39306e-315
0
11 Signal Gen~
195 171 555 0 64 64
0 11 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V4
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.89731e-315 5.34643e-315
0
7 Ground~
168 282 615 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.89731e-315 5.32571e-315
0
7 Ground~
168 282 481 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
5.89731e-315 5.30499e-315
0
11 Signal Gen~
195 171 421 0 64 64
0 14 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V3
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
5.89731e-315 5.26354e-315
0
7 Ground~
168 599 330 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
5.89731e-315 5.37752e-315
0
11 Signal Gen~
195 488 270 0 64 64
0 17 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V7
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
5.89731e-315 5.36716e-315
0
9 Inductor~
219 301 239 0 2 5
0 18 19
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
2 L2
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89731e-315 5.32571e-315
0
11 Signal Gen~
195 162 269 0 64 64
0 20 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
5.89731e-315 5.26354e-315
0
7 Ground~
168 273 329 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
5.89731e-315 0
0
9 Inductor~
219 411 88 0 2 5
0 21 22
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89731e-315 5.32571e-315
0
10 Capacitor~
219 451 125 0 2 5
0 2 22
0
0 0 848 90
8 0.9272nF
-6 0 50 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7100 0 0
2
5.89731e-315 5.30499e-315
0
7 Ground~
168 383 178 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
5.89731e-315 5.26354e-315
0
11 Signal Gen~
195 274 119 0 64 64
0 23 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400511 -1073741824 1073741824
0 814313567 814313567 939656703 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 22
20
0 16000 -2 2 0 1e-09 1e-09 3.1e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
5.89731e-315 0
0
9 Resistor~
219 573 391 0 2 5
0 8 6
0
0 0 880 0
6 3.192k
-21 -14 21 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
5.89731e-315 5.43451e-315
0
9 Resistor~
219 573 525 0 2 5
0 5 3
0
0 0 880 0
7 6.3849k
-24 -14 25 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
5.89731e-315 5.43192e-315
0
9 Resistor~
219 247 524 0 2 5
0 11 9
0
0 0 880 0
3 532
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.89731e-315 5.42933e-315
0
9 Resistor~
219 247 390 0 2 5
0 14 12
0
0 0 880 0
6 1.064k
-21 -14 21 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
5.89731e-315 5.42414e-315
0
9 Resistor~
219 564 239 0 2 5
0 17 15
0
0 0 880 0
6 2.660k
-21 -14 21 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
5.89731e-315 5.39306e-315
0
9 Resistor~
219 238 238 0 2 5
0 20 18
0
0 0 880 0
6 1.596k
-21 -14 21 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
5.89731e-315 5.38788e-315
0
9 Resistor~
219 348 87 0 2 5
0 23 21
0
0 0 880 0
6 2.128k
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
5.89731e-315 5.34643e-315
0
35
1 0 2 0 0 4096 0 14 0 0 3 2
608 610
608 606
1 2 3 0 0 8320 0 1 30 0 0 2
621 525
591 525
1 2 2 0 0 8320 0 6 15 0 0 5
676 572
676 606
537 606
537 561
528 561
2 2 4 0 0 8320 0 1 6 0 0 3
657 525
676 525
676 554
1 1 5 0 0 8320 0 15 30 0 0 4
528 551
537 551
537 525
555 525
1 0 2 0 0 0 0 13 0 0 8 2
608 476
608 472
1 2 6 0 0 8320 0 2 29 0 0 2
620 391
591 391
1 2 2 0 0 0 0 7 12 0 0 5
676 438
676 472
537 472
537 427
528 427
2 2 7 0 0 8320 0 2 7 0 0 3
656 391
676 391
676 420
1 1 8 0 0 8320 0 12 29 0 0 4
528 417
537 417
537 391
555 391
1 0 2 0 0 0 0 17 0 0 13 2
282 609
282 605
1 2 9 0 0 8320 0 4 31 0 0 3
292 523
292 524
265 524
1 2 2 0 0 0 0 9 16 0 0 5
350 572
350 605
211 605
211 560
202 560
2 2 10 0 0 8320 0 4 9 0 0 3
328 523
350 523
350 554
1 1 11 0 0 8320 0 16 31 0 0 4
202 550
211 550
211 524
229 524
1 0 2 0 0 0 0 18 0 0 18 2
282 475
282 471
1 2 12 0 0 8320 0 5 32 0 0 3
292 391
292 390
265 390
1 2 2 0 0 0 0 10 19 0 0 6
349 439
350 439
350 471
211 471
211 426
202 426
2 2 13 0 0 8320 0 5 10 0 0 4
328 391
350 391
350 421
349 421
1 1 14 0 0 8320 0 19 32 0 0 4
202 416
211 416
211 390
229 390
1 0 2 0 0 0 0 20 0 0 23 2
599 324
599 320
1 2 15 0 0 8320 0 3 33 0 0 4
610 240
609 240
609 239
582 239
1 2 2 0 0 0 0 8 21 0 0 5
667 286
667 320
528 320
528 275
519 275
2 2 16 0 0 8320 0 3 8 0 0 3
646 240
667 240
667 268
1 1 17 0 0 8320 0 21 33 0 0 4
519 265
528 265
528 239
546 239
1 0 2 0 0 0 0 24 0 0 28 2
273 323
273 319
1 2 18 0 0 8320 0 22 34 0 0 3
283 239
283 238
256 238
1 2 2 0 0 0 0 11 23 0 0 5
341 286
341 319
202 319
202 274
193 274
2 2 19 0 0 8320 0 22 11 0 0 3
319 239
341 239
341 268
1 1 20 0 0 8320 0 23 34 0 0 4
193 264
202 264
202 238
220 238
1 0 2 0 0 0 0 27 0 0 33 2
383 172
383 168
1 2 21 0 0 8320 0 25 35 0 0 3
393 88
393 87
366 87
1 2 2 0 0 0 0 26 28 0 0 6
451 134
451 168
312 168
312 123
305 123
305 124
2 2 22 0 0 8320 0 25 26 0 0 3
429 88
451 88
451 116
1 1 23 0 0 12416 0 28 35 0 0 5
305 114
305 113
312 113
312 87
330 87
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.0003125 1.25e-06 1.25e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
