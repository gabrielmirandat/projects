CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
239 130 1254 667
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.499069 0.500000
407 226 1422 494
1083744434 0
0
6 Title:
5 Name:
0
0
0
8
7 Ground~
168 268 280 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
42282.7 1
0
9 V Source~
197 323 234 0 2 5
0 3 2
0
0 0 17264 0
5 2.05V
6 0 41 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
391 0 0
2
5.89726e-315 0
0
9 V Source~
197 96 206 0 2 5
0 6 2
0
0 0 17264 0
6 3.013V
2 0 44 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3124 0 0
2
5.89726e-315 0
0
9 Resistor~
219 420 210 0 3 5
0 2 4 -1
0
0 0 880 90
4 2.2k
1 0 29 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66071556
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
5.89726e-315 0
0
9 Resistor~
219 323 188 0 2 5
0 3 4
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66070708
82 0 0 0 1 0 0 0
1 R
8157 0 0
2
5.89726e-315 0
0
9 Resistor~
219 271 160 0 2 5
0 4 5
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66069844
82 0 0 0 1 0 0 0
1 R
5572 0 0
2
5.89726e-315 0
0
9 Resistor~
219 209 214 0 3 5
0 2 5 -1
0
0 0 880 90
4 4.7k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66069048
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
5.89726e-315 0
0
9 Resistor~
219 151 160 0 2 5
0 6 5
0
0 0 880 0
3 100
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 66072404
82 0 0 0 1 0 0 0
1 R
7361 0 0
2
5.89726e-315 0
0
10
1 0 2 0 0 4096 0 1 0 0 3 2
268 274
268 260
0 2 2 0 0 4096 0 0 3 3 0 3
209 260
96 260
96 227
0 1 2 0 0 4224 0 0 7 4 0 3
323 260
209 260
209 232
2 1 2 0 0 16 0 2 4 0 0 4
323 255
323 260
420 260
420 228
1 1 3 0 0 4224 0 5 2 0 0 2
323 206
323 213
2 0 4 0 0 4096 0 5 0 0 7 2
323 170
323 160
1 2 4 0 0 4224 0 6 4 0 0 3
289 160
420 160
420 192
2 0 5 0 0 4096 0 7 0 0 9 2
209 196
209 160
2 2 5 0 0 4224 0 8 6 0 0 2
169 160
253 160
1 1 6 0 0 8320 0 3 8 0 0 3
96 185
96 160
133 160
0
0
17 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
