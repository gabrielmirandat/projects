CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
43025554 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 76 221 0 1 11
0 11
0
0 0 22368 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
1 B
-4 -30 3 -22
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.89725e-315 0
0
13 Logic Switch~
5 74 140 0 1 11
0 2
0
0 0 22368 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
1 A
-3 -30 4 -22
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3108 0 0
2
5.89725e-315 5.26354e-315
0
9 2-In AND~
219 339 41 0 3 22
0 2 3 5
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4299 0 0
2
5.89725e-315 0
0
8 2-In OR~
219 415 75 0 3 22
0 5 6 4
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9672 0 0
2
5.89725e-315 0
0
14 Logic Display~
6 913 110 0 1 2
10 15
0
0 0 56944 0
6 100MEG
-19 -24 23 -16
1 C
-4 -21 3 -13
1 C
-4 -41 3 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 1 0 0
1 L
7876 0 0
2
5.89725e-315 5.30499e-315
0
14 Logic Display~
6 657 206 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89725e-315 5.32571e-315
0
14 Logic Display~
6 654 54 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89725e-315 5.34643e-315
0
8 2-In OR~
219 487 114 0 3 22
0 4 14 3
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7100 0 0
2
5.89725e-315 5.3568e-315
0
8 2-In OR~
219 490 272 0 3 22
0 7 8 13
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3820 0 0
2
5.89725e-315 5.36716e-315
0
8 2-In OR~
219 409 227 0 3 22
0 10 9 7
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7678 0 0
2
5.89725e-315 5.37752e-315
0
9 Inverter~
13 590 245 0 2 22
0 13 16
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
961 0 0
2
5.89725e-315 5.38788e-315
0
9 Inverter~
13 173 94 0 2 22
0 2 12
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3178 0 0
2
5.89725e-315 5.39306e-315
0
9 2-In AND~
219 857 158 0 3 22
0 3 16 15
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3409 0 0
2
5.89725e-315 5.39824e-315
0
9 2-In AND~
219 342 205 0 3 22
0 12 13 10
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
5.89725e-315 5.40342e-315
0
9 2-In AND~
219 342 313 0 3 22
0 12 11 8
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8885 0 0
2
5.89725e-315 5.4086e-315
0
9 2-In AND~
219 342 258 0 3 22
0 11 13 9
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3780 0 0
2
5.89725e-315 5.41378e-315
0
9 2-In AND~
219 341 149 0 3 22
0 2 11 14
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9265 0 0
2
5.89725e-315 5.41896e-315
0
9 2-In AND~
219 341 94 0 3 22
0 11 3 6
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9442 0 0
2
5.89725e-315 5.42414e-315
0
27
0 1 2 0 0 8192 0 0 3 6 0 3
129 95
129 32
315 32
0 2 3 0 0 4096 0 0 3 21 0 3
274 104
274 50
315 50
3 1 4 0 0 8320 0 4 8 0 0 4
448 75
463 75
463 105
474 105
1 3 5 0 0 4224 0 4 3 0 0 4
402 66
375 66
375 41
360 41
3 2 6 0 0 12416 0 18 4 0 0 4
362 94
375 94
375 84
402 84
0 1 2 0 0 0 0 0 12 7 0 3
129 140
129 94
158 94
1 1 2 0 0 4224 0 2 17 0 0 2
86 140
317 140
3 1 7 0 0 8320 0 10 9 0 0 4
442 227
454 227
454 263
477 263
3 2 8 0 0 12416 0 15 9 0 0 4
363 313
375 313
375 281
477 281
3 2 9 0 0 8320 0 16 10 0 0 4
363 258
375 258
375 236
396 236
3 1 10 0 0 12416 0 14 10 0 0 4
363 205
375 205
375 218
396 218
0 2 11 0 0 8192 0 0 15 14 0 3
222 249
222 322
318 322
0 1 12 0 0 8320 0 0 15 15 0 3
204 196
204 304
318 304
0 1 11 0 0 0 0 0 16 20 0 3
222 221
222 249
318 249
2 1 12 0 0 0 0 12 14 0 0 4
194 94
204 94
204 196
318 196
2 0 13 0 0 4096 0 16 0 0 17 2
318 267
247 267
0 2 13 0 0 8320 0 0 14 25 0 5
556 272
556 384
247 384
247 214
318 214
3 2 14 0 0 12416 0 17 8 0 0 4
362 149
375 149
375 123
474 123
2 0 11 0 0 0 0 17 0 0 20 2
317 158
222 158
1 1 11 0 0 8320 0 18 1 0 0 4
317 85
222 85
222 221
88 221
0 2 3 0 0 8320 0 0 18 23 0 5
699 114
699 359
274 359
274 103
317 103
3 1 15 0 0 4224 0 13 5 0 0 3
878 158
913 158
913 128
0 1 3 0 0 0 0 0 13 27 0 4
653 114
806 114
806 149
833 149
2 2 16 0 0 4224 0 11 13 0 0 4
611 245
806 245
806 167
833 167
0 1 13 0 0 0 0 0 11 26 0 3
556 272
556 245
575 245
3 1 13 0 0 0 0 9 6 0 0 3
523 272
657 272
657 224
3 1 3 0 0 0 0 8 7 0 0 3
520 114
654 114
654 72
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
