CircuitMaker Text
5.6
Probes: 1
L1_2
Transient Analysis
0 419 204 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 170 30 280 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
98 C:\Users\Marina\Desktop\Backup\4� semestre\Sistemas digitais 1\Laborat�rio\CircuitMakerfim\BOM.DAT
0 7
2 4 0.500000 0.500000
176 79 1364 393
1083966130 0
0
6 Title:
5 Name:
0
0
0
10
5 SAVE-
218 309 202 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
47 0 0
2
42127.9 0
0
5 SCOPE
12 157 192 0 1 11
0 3
0
0 0 57584 0
2 A2
-8 -4 6 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5391 0 0
2
42127.6 0
0
5 SCOPE
12 282 191 0 1 11
0 4
0
0 0 57584 0
2 A1
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3945 0 0
2
42127.6 0
0
5 SCOPE
12 381 190 0 1 11
0 5
0
0 0 57584 0
1 A
-4 -4 3 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5628 0 0
2
42127.6 0
0
9 Inductor~
219 381 237 0 2 5
0 2 5
0
0 0 848 602
2 6H
9 -4 23 4
2 L2
10 -14 24 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
3283 0 0
2
42127.6 0
0
9 Inductor~
219 338 203 0 2 5
0 4 5
0
0 0 848 0
5 470uH
-18 -17 17 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
7481 0 0
2
42127.6 0
0
7 Ground~
168 262 285 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
339 0 0
2
42127.6 0
0
11 Signal Gen~
195 124 245 0 19 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1067785912 1114636288 0 1067819467
20
1.29 60 0 1.294 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -1.29/1.29V
-39 -30 38 -22
2 V1
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 1.294 60 0 0) AC 1.29 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 1 0 0
1 V
3593 0 0
2
42127.6 0
0
9 Resistor~
219 451 235 0 3 5
0 2 5 -1
0
0 0 880 90
6 5.051k
-6 0 36 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4568 0 0
2
42127.6 0
0
9 Resistor~
219 236 202 0 2 5
0 3 4
0
0 0 880 0
6 1.051k
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3338 0 0
2
42127.6 0
0
11
1 0 3 0 0 4096 0 2 0 0 5 2
157 204
155 204
1 0 4 0 0 4096 0 3 0 0 8 2
282 203
282 202
1 0 5 0 0 4096 0 4 0 0 6 2
381 202
381 203
1 0 2 0 0 4096 0 7 0 0 10 2
262 279
262 280
1 1 3 0 0 8320 0 8 10 0 0 3
155 240
155 202
218 202
2 0 5 0 0 4096 0 5 0 0 11 2
381 219
381 203
2 0 5 0 0 0 0 9 0 0 11 2
451 217
451 209
1 2 4 0 0 8320 0 6 10 0 0 3
320 203
320 202
254 202
1 0 2 0 0 4096 0 5 0 0 10 2
381 255
381 280
1 2 2 0 0 8320 0 9 8 0 0 4
451 253
451 280
155 280
155 250
2 2 5 0 0 4224 0 6 9 0 0 3
356 203
451 203
451 217
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.0833333 0.000333333 0.000333333
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
