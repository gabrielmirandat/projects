CircuitMaker Text
5.6
Probes: 3
R15_2
Transient Analysis
0 1023 176 16512
R15_1
Transient Analysis
1 963 144 16711935
R17_1
Transient Analysis
2 966 209 255
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 40 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
56
7 Ground~
168 347 428 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
449 0 0
2
42334.5 0
0
11 Signal Gen~
195 195 224 0 64 64
0 5 7 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1073741824 0 1084227584
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 2 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -5/5V
-18 -30 17 -22
3 V11
-10 -40 11 -32
0
0
35 %D %1 %2 DC 0 SIN(0 5 2 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8761 0 0
2
5.89732e-315 0
0
11 Signal Gen~
195 189 124 0 64 64
0 6 5 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1073741824 0 1084227584
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 2 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -5/5V
-18 -30 17 -22
3 V10
-10 -40 11 -32
0
0
35 %D %1 %2 DC 0 SIN(0 5 2 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6748 0 0
2
5.89732e-315 0
0
11 Signal Gen~
195 107 286 0 19 64
0 5 8 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1073741824 0 1084227584
20
1 2 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -5/5V
-18 -30 17 -22
2 V9
-7 -40 7 -32
0
0
35 %D %1 %2 DC 0 SIN(0 5 2 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7393 0 0
2
5.89732e-315 0
0
5 SCOPE
12 1117 147 0 1 11
0 9
0
0 0 57584 0
5 SA�DA
-18 -4 17 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7699 0 0
2
5.89732e-315 0
0
10 Capacitor~
219 324 67 0 2 5
0 24 21
0
0 0 336 0
4 47nF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6638 0 0
2
5.89732e-315 5.37752e-315
0
10 Capacitor~
219 322 217 0 2 5
0 23 20
0
0 0 336 0
4 47nF
-14 -18 14 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4595 0 0
2
5.89732e-315 5.36716e-315
0
10 Capacitor~
219 430 145 0 2 5
0 2 22
0
0 0 336 90
4 33pF
-43 -3 -15 5
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9395 0 0
2
5.89732e-315 5.3568e-315
0
10 Capacitor~
219 453 157 0 2 5
0 4 2
0
0 0 336 180
4 33pF
-14 -18 14 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3303 0 0
2
5.89732e-315 5.34643e-315
0
10 Capacitor~
219 580 168 0 2 5
0 3 15
0
0 0 336 90
5 330pF
9 -5 44 3
2 C5
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4498 0 0
2
5.89732e-315 5.32571e-315
0
10 Capacitor~
219 652 155 0 2 5
0 2 3
0
0 0 336 180
4 33pF
-14 -18 14 -10
2 C6
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9728 0 0
2
5.89732e-315 5.30499e-315
0
10 Capacitor~
219 675 139 0 2 5
0 2 15
0
0 0 336 90
4 33pF
12 -5 40 3
2 C7
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3789 0 0
2
5.89732e-315 5.26354e-315
0
6 Diode~
219 835 228 0 2 5
0 19 18
0
0 0 80 270
5 DIODE
-18 -18 17 -10
2 D4
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3978 0 0
2
5.89732e-315 5.26354e-315
0
6 Diode~
219 812 229 0 2 5
0 18 19
0
0 0 80 90
5 DIODE
-18 -18 17 -10
2 D3
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3494 0 0
2
5.89732e-315 0
0
6 Diode~
219 831 100 0 2 5
0 17 16
0
0 0 80 270
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3507 0 0
2
5.89732e-315 5.26354e-315
0
6 Diode~
219 808 101 0 2 5
0 16 17
0
0 0 80 90
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
5151 0 0
2
5.89732e-315 0
0
10 Op-Amp5:A~
219 872 88 0 5 11
0 17 16 27 28 10
0
0 0 80 0
5 TL064
15 -25 50 -17
2 U3
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3701 0 0
2
5.89732e-315 5.30499e-315
0
2 +V
167 873 114 0 1 3
0 28
0
0 0 53616 180
4 -15V
3 -7 31 1
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8585 0 0
2
5.89732e-315 5.26354e-315
0
2 +V
167 872 67 0 1 3
0 27
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8809 0 0
2
5.89732e-315 0
0
2 +V
167 876 224 0 1 3
0 29
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5993 0 0
2
5.89732e-315 0
0
2 +V
167 987 155 0 1 3
0 30
0
0 0 53616 0
3 15V
-11 -22 10 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8654 0 0
2
5.89732e-315 0
0
2 +V
167 987 201 0 1 3
0 31
0
0 0 53616 180
4 -15V
3 -7 31 1
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7223 0 0
2
5.89732e-315 0
0
2 +V
167 875 268 0 1 3
0 32
0
0 0 53616 180
4 -15V
3 -7 31 1
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3641 0 0
2
5.89732e-315 0
0
8 Op-Amp5~
219 986 175 0 5 11
0 26 25 30 31 9
0
0 0 80 0
5 TL064
15 -25 50 -17
3 U4B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP14
26

0 5 6 4 11 7 3 2 4 11
1 5 6 4 11 7 10 9 4 11
8 12 13 4 11 14 0
88 0 0 0 4 2 1 0
1 U
3104 0 0
2
5.89732e-315 0
0
8 Op-Amp5~
219 875 243 0 5 11
0 18 19 29 32 12
0
0 0 80 0
5 TL064
15 -25 50 -17
3 U4A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP14
26

0 3 2 4 11 1 3 2 4 11
1 5 6 4 11 7 10 9 4 11
8 12 13 4 11 14 62
88 0 0 0 4 1 1 0
1 U
3296 0 0
2
5.89732e-315 0
0
10 Op-Amp5:A~
219 648 357 0 5 11
0 38 35 37 2 36
0
0 0 80 180
5 TL064
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 512 1 0 0 0
1 U
8534 0 0
2
5.89732e-315 5.38788e-315
0
2 +V
167 648 395 0 1 3
0 37
0
0 0 53616 180
3 15V
6 -7 27 1
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
949 0 0
2
5.89732e-315 5.3568e-315
0
2 +V
167 768 389 0 1 3
0 34
0
0 0 53616 180
3 15V
6 -7 27 1
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3371 0 0
2
5.89732e-315 5.32571e-315
0
10 Op-Amp5:A~
219 768 350 0 5 11
0 11 33 34 2 33
0
0 0 80 180
5 TL064
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
7311 0 0
2
5.89732e-315 5.26354e-315
0
9 Resistor~
219 1045 311 0 2 5
0 11 10
0
0 0 368 90
3 10k
7 -5 28 3
3 R27
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.89732e-315 0
0
9 Resistor~
219 863 316 0 2 5
0 11 12
0
0 0 368 90
3 10k
7 -5 28 3
3 R26
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3526 0 0
2
5.89732e-315 0
0
9 Resistor~
219 726 164 0 2 5
0 13 14
0
0 0 368 90
2 4k
8 -5 22 3
3 R25
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4129 0 0
2
5.89732e-315 0
0
9 Resistor~
219 762 246 0 2 5
0 3 18
0
0 0 368 0
2 1k
-7 -14 7 -6
3 R24
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6278 0 0
2
5.89732e-315 0
0
9 Resistor~
219 763 215 0 2 5
0 13 19
0
0 0 368 0
2 1k
-7 -14 7 -6
3 R23
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3482 0 0
2
5.89732e-315 0
0
9 Resistor~
219 761 120 0 2 5
0 14 16
0
0 0 368 0
2 1k
-7 -14 7 -6
3 R22
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8323 0 0
2
5.89732e-315 0
0
9 Resistor~
219 757 76 0 2 5
0 15 17
0
0 0 368 0
2 1k
-7 -14 7 -6
3 R21
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3984 0 0
2
5.89732e-315 0
0
9 Resistor~
219 262 96 0 2 5
0 6 24
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7622 0 0
2
5.89732e-315 5.42414e-315
0
9 Resistor~
219 324 134 0 2 5
0 24 21
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
816 0 0
2
5.89732e-315 5.41896e-315
0
9 Resistor~
219 324 282 0 2 5
0 23 20
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4656 0 0
2
5.89732e-315 5.41378e-315
0
9 Resistor~
219 261 254 0 2 5
0 7 23
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6356 0 0
2
5.89732e-315 5.4086e-315
0
9 Resistor~
219 386 117 0 2 5
0 21 22
0
0 0 368 0
5 63.4k
-17 -14 18 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7479 0 0
2
5.89732e-315 5.40342e-315
0
9 Resistor~
219 500 116 0 2 5
0 22 15
0
0 0 368 0
5 63.4k
-17 -14 18 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5690 0 0
2
5.89732e-315 5.39824e-315
0
9 Resistor~
219 436 243 0 2 5
0 20 4
0
0 0 368 0
5 63.4k
-17 -14 18 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5617 0 0
2
5.89732e-315 5.39306e-315
0
9 Resistor~
219 517 243 0 2 5
0 4 3
0
0 0 368 0
5 63.4k
-17 -14 18 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3903 0 0
2
5.89732e-315 5.38788e-315
0
9 Resistor~
219 886 190 0 2 5
0 13 12
0
0 0 368 0
3 20k
-10 -14 11 -6
3 R20
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4452 0 0
2
5.89732e-315 0
0
9 Resistor~
219 880 154 0 2 5
0 14 10
0
0 0 368 0
3 20k
-10 -14 11 -6
3 R19
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6282 0 0
2
5.89732e-315 0
0
9 Resistor~
219 938 254 0 2 5
0 12 26
0
0 0 368 0
3 10k
-10 -14 11 -6
3 R18
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7187 0 0
2
5.89732e-315 0
0
9 Resistor~
219 979 254 0 4 5
0 26 2 0 -1
0
0 0 368 0
3 10k
-10 -14 11 -6
3 R17
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6866 0 0
2
5.89732e-315 0
0
9 Resistor~
219 950 107 0 2 5
0 10 25
0
0 0 368 0
3 10k
-10 -14 11 -6
3 R16
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7670 0 0
2
5.89732e-315 0
0
9 Resistor~
219 1000 106 0 2 5
0 25 9
0
0 0 368 0
3 10k
-10 -14 11 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
951 0 0
2
5.89732e-315 0
0
9 Resistor~
219 586 345 0 2 5
0 8 36
0
0 0 368 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9536 0 0
2
5.89732e-315 5.41896e-315
0
9 Resistor~
219 610 394 0 3 5
0 2 36 -1
0
0 0 368 90
2 1M
8 -5 22 3
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5495 0 0
2
5.89732e-315 5.41378e-315
0
9 Resistor~
219 649 303 0 2 5
0 36 35
0
0 0 368 0
2 1M
-7 -14 7 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8152 0 0
2
5.89732e-315 5.4086e-315
0
9 Resistor~
219 725 351 0 2 5
0 35 33
0
0 0 368 0
3 10k
-10 -14 11 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6223 0 0
2
5.89732e-315 5.40342e-315
0
9 Resistor~
219 746 405 0 3 5
0 2 33 -1
0
0 0 368 90
2 1M
8 -5 22 3
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5441 0 0
2
5.89732e-315 5.39824e-315
0
9 Resistor~
219 818 397 0 3 5
0 2 11 -1
0
0 0 368 90
2 1M
8 -5 22 3
3 R14
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3189 0 0
2
5.89732e-315 5.39306e-315
0
82
0 0 3 0 0 4096 0 0 0 2 3 2
614 181
614 246
1 2 3 0 0 0 0 10 11 0 0 5
580 177
580 181
635 181
635 155
643 155
1 2 3 0 0 4224 0 33 44 0 0 4
744 246
543 246
543 243
535 243
0 0 2 0 0 4096 0 0 0 13 5 3
710 423
710 155
675 155
1 1 2 0 0 0 0 12 11 0 0 3
675 148
675 155
661 155
0 0 2 0 0 0 0 0 0 8 14 3
430 157
374 157
374 412
1 0 4 0 0 8320 0 9 0 0 46 3
462 157
474 157
474 244
1 2 2 0 0 0 0 8 9 0 0 3
430 154
430 157
444 157
2 0 2 0 0 0 0 48 0 0 12 3
997 254
997 434
818 434
4 0 2 0 0 0 0 29 0 0 11 3
768 337
768 316
648 316
4 0 2 0 0 0 0 26 0 0 14 4
648 344
648 315
517 315
517 412
1 0 2 0 0 8320 0 56 0 0 14 4
818 415
818 434
527 434
527 412
1 0 2 0 0 0 0 55 0 0 14 3
746 423
533 423
533 412
1 1 2 0 0 0 0 1 52 0 0 3
347 422
347 412
610 412
1 0 5 0 0 4224 0 4 0 0 18 3
138 281
138 176
241 176
1 1 6 0 0 8320 0 3 37 0 0 4
220 119
236 119
236 96
244 96
2 1 7 0 0 8320 0 2 40 0 0 4
226 229
235 229
235 254
243 254
1 2 5 0 0 0 0 2 3 0 0 4
226 219
241 219
241 129
220 129
2 1 8 0 0 4224 0 4 51 0 0 4
138 291
560 291
560 345
568 345
0 1 9 0 0 4224 0 0 5 59 0 3
1026 175
1117 175
1117 159
2 0 10 0 0 4224 0 30 0 0 57 4
1045 293
1045 72
902 72
902 107
0 1 11 0 0 4224 0 0 30 24 0 3
863 356
1045 356
1045 329
2 0 12 0 0 4096 0 31 0 0 55 3
863 298
913 298
913 254
0 1 11 0 0 0 0 0 31 70 0 3
818 356
863 356
863 334
1 0 13 0 0 4224 0 45 0 0 26 2
868 190
725 190
1 1 13 0 0 0 0 34 32 0 0 5
745 215
725 215
725 190
726 190
726 182
1 0 14 0 0 8320 0 46 0 0 28 5
862 154
862 127
733 127
733 126
725 126
1 2 14 0 0 0 0 35 32 0 0 5
743 120
725 120
725 126
726 126
726 146
1 0 15 0 0 4224 0 36 0 0 44 3
739 76
627 76
627 117
0 2 16 0 0 12288 0 0 17 37 0 5
830 118
830 114
846 114
846 94
854 94
0 1 17 0 0 4096 0 0 17 36 0 2
831 82
854 82
0 1 18 0 0 8192 0 0 25 38 0 3
833 251
833 249
857 249
0 2 19 0 0 12288 0 0 25 41 0 5
835 210
835 214
849 214
849 237
857 237
2 0 17 0 0 4224 0 36 0 0 36 4
775 76
803 76
803 82
808 82
2 0 16 0 0 4224 0 35 0 0 37 3
779 120
811 120
811 118
2 1 17 0 0 0 0 16 15 0 0 4
808 91
808 82
831 82
831 90
1 2 16 0 0 0 0 16 15 0 0 4
808 111
808 118
831 118
831 110
1 2 18 0 0 0 0 14 13 0 0 4
812 239
812 251
835 251
835 238
2 1 18 0 0 4224 0 33 14 0 0 3
780 246
812 246
812 239
2 0 19 0 0 4224 0 34 0 0 41 2
781 215
812 215
2 1 19 0 0 0 0 14 13 0 0 4
812 219
812 210
835 210
835 218
1 0 20 0 0 4224 0 43 0 0 49 2
418 243
345 243
1 0 21 0 0 4224 0 41 0 0 52 2
368 117
346 117
2 0 15 0 0 0 0 12 0 0 45 3
675 130
675 117
579 117
2 2 15 0 0 0 0 10 42 0 0 5
580 159
580 117
579 117
579 116
518 116
2 1 4 0 0 128 0 43 44 0 0 5
454 243
454 244
474 244
474 243
499 243
0 2 22 0 0 4096 0 0 8 48 0 2
430 117
430 136
2 1 22 0 0 12416 0 41 42 0 0 4
404 117
430 117
430 116
482 116
2 2 20 0 0 0 0 7 39 0 0 4
331 217
345 217
345 282
342 282
0 1 23 0 0 4224 0 0 39 51 0 3
294 217
294 282
306 282
2 1 23 0 0 0 0 40 7 0 0 4
279 254
294 254
294 217
313 217
2 2 21 0 0 8320 0 6 38 0 0 4
333 67
346 67
346 134
342 134
0 1 24 0 0 4224 0 0 38 54 0 3
295 96
295 134
306 134
2 1 24 0 0 0 0 37 6 0 0 4
280 96
295 96
295 67
315 67
2 0 12 0 0 8320 0 45 0 0 56 3
904 190
913 190
913 254
1 5 12 0 0 0 0 47 25 0 0 4
920 254
901 254
901 243
893 243
2 0 10 0 0 0 0 46 0 0 58 3
898 154
902 154
902 107
1 5 10 0 0 0 0 49 17 0 0 4
932 107
898 107
898 88
890 88
5 2 9 0 0 0 0 24 50 0 0 4
1004 175
1026 175
1026 106
1018 106
1 0 25 0 0 4096 0 50 0 0 63 3
982 106
973 106
973 107
1 0 26 0 0 4096 0 48 0 0 62 2
961 254
962 254
1 2 26 0 0 8320 0 24 47 0 0 6
968 181
964 181
964 248
962 248
962 254
956 254
2 2 25 0 0 8320 0 24 49 0 0 6
968 169
964 169
964 115
973 115
973 107
968 107
1 3 27 0 0 4224 0 19 17 0 0 2
872 76
872 75
1 4 28 0 0 4224 0 18 17 0 0 3
873 99
873 101
872 101
1 3 29 0 0 4224 0 20 25 0 0 3
876 233
876 230
875 230
1 3 30 0 0 4224 0 21 24 0 0 3
987 164
987 162
986 162
1 4 31 0 0 4224 0 22 24 0 0 3
987 186
987 188
986 188
1 4 32 0 0 4224 0 23 25 0 0 2
875 253
875 256
1 2 11 0 0 0 0 29 56 0 0 3
786 356
818 356
818 379
1 0 2 0 0 0 0 56 0 0 0 4
818 415
818 417
817 417
817 416
2 2 33 0 0 8320 0 29 54 0 0 4
786 344
786 309
743 309
743 351
1 3 34 0 0 4224 0 28 29 0 0 2
768 374
768 363
1 0 2 0 0 0 0 55 0 0 0 4
746 423
746 425
745 425
745 424
2 0 33 0 0 0 0 55 0 0 76 2
746 387
746 351
5 2 33 0 0 0 0 29 54 0 0 6
750 350
746 350
746 351
742 351
742 351
743 351
1 0 35 0 0 4096 0 54 0 0 78 2
707 351
680 351
2 2 35 0 0 8320 0 26 53 0 0 4
666 351
680 351
680 303
667 303
5 0 36 0 0 4096 0 26 0 0 81 2
630 357
610 357
2 0 36 0 0 0 0 51 0 0 81 2
604 345
610 345
2 1 36 0 0 4224 0 52 53 0 0 3
610 376
610 303
631 303
1 3 37 0 0 4224 0 27 26 0 0 2
648 380
648 370
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 2.5 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
