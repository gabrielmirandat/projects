CircuitMaker Text
5.6
Probes: 6
V1_1
Transient Analysis
0 327 71 65280
L_1
Transient Analysis
1 373 73 65535
L_2
Transient Analysis
2 442 72 16776960
V1_1
Operating Point
0 328 75 65280
L_1
Operating Point
1 376 74 65535
L_2
Operating Point
2 438 72 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 79 1364 384
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
25
9 Inductor~
219 579 300 0 2 5
0 3 4
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
2 L4
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
5130 0 0
2
5.89732e-315 5.34643e-315
0
10 Capacitor~
219 619 337 0 2 5
0 2 4
0
0 0 848 90
8 0.9272nF
-6 0 50 8
2 C4
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
391 0 0
2
5.89732e-315 5.32571e-315
0
7 Ground~
168 551 390 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.89732e-315 5.30499e-315
0
11 Signal Gen~
195 442 331 0 64 64
0 5 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1218282720 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2255372
20
0 322599 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V5
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 500m 322.6k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3421 0 0
2
5.89732e-315 5.26354e-315
0
9 Inductor~
219 576 186 0 2 5
0 6 7
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
2 L3
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89732e-315 5.34643e-315
0
10 Capacitor~
219 616 223 0 2 5
0 2 7
0
0 0 848 90
8 0.9272nF
-6 0 50 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5572 0 0
2
5.89732e-315 5.32571e-315
0
7 Ground~
168 548 276 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.89732e-315 5.30499e-315
0
11 Signal Gen~
195 439 217 0 64 64
0 8 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1215055616 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 241948 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V4
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 500m 241.9k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89732e-315 5.26354e-315
0
9 Inductor~
219 248 308 0 2 5
0 9 10
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
2 L2
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89732e-315 5.32571e-315
0
10 Capacitor~
219 288 345 0 2 5
0 2 10
0
0 0 848 90
8 0.9272nF
-6 0 50 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
972 0 0
2
5.89732e-315 5.30499e-315
0
7 Ground~
168 220 398 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
5.89732e-315 5.26354e-315
0
11 Signal Gen~
195 111 339 0 64 64
0 11 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1201505536 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 80650 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 500m 80.65k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.89732e-315 0
0
9 Inductor~
219 250 187 0 2 5
0 12 13
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.89732e-315 5.34643e-315
0
10 Capacitor~
219 290 224 0 2 5
0 2 13
0
0 0 848 90
8 0.9272nF
-6 0 50 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4597 0 0
2
5.89732e-315 5.32571e-315
0
7 Ground~
168 222 277 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
5.89732e-315 5.30499e-315
0
11 Signal Gen~
195 113 218 0 64 64
0 14 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1193116928 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 40325 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 500m 40.33k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.89732e-315 5.26354e-315
0
11 Signal Gen~
195 276 105 0 64 64
0 17 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1209894144 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 161300 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 500m 161.3k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
5.89732e-315 5.32571e-315
0
7 Ground~
168 385 164 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
5.89732e-315 5.30499e-315
0
10 Capacitor~
219 453 111 0 2 5
0 2 16
0
0 0 848 90
8 0.9272nF
-6 0 50 8
1 C
18 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
317 0 0
2
5.89732e-315 5.26354e-315
0
9 Inductor~
219 413 74 0 2 5
0 15 16
0
0 0 848 0
6 1.05mH
-21 -17 21 -9
1 L
-4 -27 3 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89732e-315 0
0
9 Resistor~
219 516 299 0 2 5
0 5 3
0
0 0 880 0
6 2.128k
-21 -14 21 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4299 0 0
2
5.89732e-315 0
0
9 Resistor~
219 513 185 0 2 5
0 8 6
0
0 0 880 0
6 2.128k
-21 -14 21 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
5.89732e-315 0
0
9 Resistor~
219 185 307 0 2 5
0 11 9
0
0 0 880 0
6 2.128k
-21 -14 21 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
5.89732e-315 0
0
9 Resistor~
219 187 186 0 2 5
0 14 12
0
0 0 880 0
6 2.128k
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
5.89732e-315 0
0
9 Resistor~
219 350 73 0 2 5
0 17 15
0
0 0 880 0
6 2.128k
-21 -14 21 -6
1 R
-4 -24 3 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
5.89732e-315 5.34643e-315
0
25
1 0 2 0 0 4096 0 3 0 0 3 2
551 384
551 380
1 2 3 0 0 8320 0 1 21 0 0 3
561 300
561 299
534 299
1 2 2 0 0 8320 0 2 4 0 0 6
619 346
619 380
480 380
480 335
473 335
473 336
2 2 4 0 0 8320 0 1 2 0 0 3
597 300
619 300
619 328
1 1 5 0 0 12416 0 4 21 0 0 5
473 326
473 325
480 325
480 299
498 299
1 0 2 0 0 0 0 7 0 0 8 2
548 270
548 266
1 2 6 0 0 8320 0 5 22 0 0 3
558 186
558 185
531 185
1 2 2 0 0 0 0 6 8 0 0 6
616 232
616 266
477 266
477 221
470 221
470 222
2 2 7 0 0 8320 0 5 6 0 0 3
594 186
616 186
616 214
1 1 8 0 0 12416 0 8 22 0 0 5
470 212
470 211
477 211
477 185
495 185
1 0 2 0 0 0 0 11 0 0 13 2
220 392
220 388
1 2 9 0 0 8320 0 9 23 0 0 3
230 308
230 307
203 307
1 2 2 0 0 0 0 10 12 0 0 6
288 354
288 388
149 388
149 343
142 343
142 344
2 2 10 0 0 8320 0 9 10 0 0 3
266 308
288 308
288 336
1 1 11 0 0 12416 0 12 23 0 0 5
142 334
142 333
149 333
149 307
167 307
1 0 2 0 0 0 0 15 0 0 18 2
222 271
222 267
1 2 12 0 0 8320 0 13 24 0 0 3
232 187
232 186
205 186
1 2 2 0 0 0 0 14 16 0 0 6
290 233
290 267
151 267
151 222
144 222
144 223
2 2 13 0 0 8320 0 13 14 0 0 3
268 187
290 187
290 215
1 1 14 0 0 12416 0 16 24 0 0 5
144 213
144 212
151 212
151 186
169 186
1 0 2 0 0 0 0 18 0 0 23 2
385 158
385 154
1 2 15 0 0 8320 0 20 25 0 0 3
395 74
395 73
368 73
1 2 2 0 0 0 0 19 17 0 0 6
453 120
453 154
314 154
314 109
307 109
307 110
2 2 16 0 0 8320 0 20 19 0 0 3
431 74
453 74
453 102
1 1 17 0 0 12416 0 17 25 0 0 5
307 100
307 99
314 99
314 73
332 73
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.000123993 2.47985e-07 2.47985e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
