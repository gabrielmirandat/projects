CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 70 10
341 118 1356 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
509 214 622 311
43024562 0
0
6 Title:
5 Name:
0
0
0
54
13 Logic Switch~
5 175 399 0 1 11
0 21
0
0 0 21344 0
2 0V
-5 -16 9 -8
2 T1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89727e-315 0
0
13 Logic Switch~
5 107 99 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
3 LEU
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89727e-315 5.39824e-315
0
13 Logic Switch~
5 103 136 0 1 11
0 34
0
0 0 21344 0
2 0V
-5 -16 9 -8
2 SO
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89727e-315 5.39306e-315
0
13 Logic Switch~
5 105 212 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
3 SOK
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89727e-315 5.38788e-315
0
13 Logic Switch~
5 102 176 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
3 TOK
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89727e-315 5.37752e-315
0
13 Logic Switch~
5 103 325 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
1 T
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89727e-315 5.36716e-315
0
13 Logic Switch~
5 104 288 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
2 HP
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89727e-315 5.3568e-315
0
13 Logic Switch~
5 103 249 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-5 -16 9 -8
3 MOK
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.89727e-315 5.34643e-315
0
8 2-In OR~
219 931 133 0 3 22
0 4 5 3
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U12C
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
4747 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 1373 65 0 1 2
10 12
0
0 0 53872 0
6 100MEG
-199 -55 -157 -47
2 LT
-5 -21 9 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89727e-315 5.26354e-315
0
14 Logic Display~
6 1425 62 0 1 2
10 11
0
0 0 53872 0
6 100MEG
-22 -36 20 -28
2 LS
-5 -21 9 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89727e-315 0
0
9 Inverter~
13 1160 284 0 2 22
0 10 11
0
0 0 608 0
6 74LS04
16 -24 58 -16
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
9998 0 0
2
5.89727e-315 0
0
9 Inverter~
13 1159 213 0 2 22
0 8 13
0
0 0 608 0
6 74LS04
18 -27 60 -19
4 U14B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
3536 0 0
2
5.89727e-315 5.26354e-315
0
9 Inverter~
13 1160 248 0 2 22
0 9 12
0
0 0 608 0
6 74LS04
9 -26 51 -18
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
4597 0 0
2
5.89727e-315 0
0
9 Inverter~
13 1159 180 0 2 22
0 7 14
0
0 0 608 0
6 74LS04
6 -28 48 -20
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3835 0 0
2
5.89727e-315 0
0
9 Inverter~
13 1158 144 0 2 22
0 6 15
0
0 0 608 0
6 74LS04
8 -29 50 -21
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3670 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 1331 65 0 1 2
10 13
0
0 0 53872 0
6 100MEG
16 -34 58 -26
3 LER
-9 -21 12 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 1288 67 0 1 2
10 14
0
0 0 53872 0
6 100MEG
15 -50 57 -42
3 AVG
-9 -21 12 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 1244 64 0 1 2
10 15
0
0 0 53872 0
6 100MEG
23 -35 65 -27
4 RETR
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89727e-315 0
0
7 Ground~
168 997 112 0 1 3
0 2
0
0 0 53344 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
5.89727e-315 0
0
8 2-In OR~
219 948 206 0 3 22
0 18 17 5
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U12B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
4299 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 1204 64 0 1 2
10 3
0
0 0 53872 0
6 100MEG
12 -37 54 -29
4 LDHD
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89727e-315 0
0
14 Logic Display~
6 1166 64 0 1 2
10 3
0
0 0 53872 0
6 100MEG
-34 -40 8 -32
2 MT
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89727e-315 0
0
2 +V
167 254 523 0 1 3
0 22
0
0 0 54240 180
3 10V
6 -2 27 6
2 V4
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6369 0 0
2
5.89727e-315 0
0
2 +V
167 254 388 0 1 3
0 23
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9172 0 0
2
5.89727e-315 0
0
5 7474~
219 254 474 0 6 22
0 23 21 20 22 49 19
0
0 0 4704 0
4 7474
7 -60 35 -52
4 U13A
7 -71 35 -63
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 9 0
1 U
7100 0 0
2
5.89727e-315 0
0
7 Pulser~
4 156 456 0 10 12
0 50 51 52 20 0 0 10 10 2
8
0
0 0 4640 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3820 0 0
2
5.89727e-315 0
0
2 +V
167 659 233 0 1 3
0 24
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
5.89727e-315 0
0
7 Ground~
168 739 309 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
5.89727e-315 0
0
8 2-In OR~
219 547 512 0 3 22
0 28 27 26
0
0 0 608 0
6 74LS32
18 -34 60 -26
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3178 0 0
2
5.89727e-315 0
0
9 Inverter~
13 330 305 0 2 22
0 27 33
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U5D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3409 0 0
2
5.89727e-315 0
0
7 74LS151
20 259 148 0 14 29
0 53 54 36 34 37 38 39 40 2
4 17 18 28 55
0
0 0 4832 0
7 74LS151
-24 -70 25 -62
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3951 0 0
2
5.89727e-315 5.32571e-315
0
7 74LS153
119 258 303 0 14 29
0 35 34 56 57 17 18 58 59 60
61 2 62 27 63
0
0 0 4832 0
7 74LS153
-24 -70 25 -62
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
8885 0 0
2
5.89727e-315 5.30499e-315
0
7 Ground~
168 334 85 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3780 0 0
2
5.89727e-315 5.26354e-315
0
7 Ground~
168 331 231 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
5.89727e-315 0
0
7 74LS194
49 738 217 0 14 29
0 19 30 29 2 26 24 2 2 25
2 18 17 4 16
0
0 0 4832 0
7 74LS194
-40 -69 9 -61
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9442 0 0
2
5.89727e-315 5.43192e-315
0
14 Logic Display~
6 890 85 0 1 2
10 18
0
0 0 53872 0
6 100MEG
14 -13 56 -5
2 QA
-8 -29 6 -21
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89727e-315 5.42933e-315
0
14 Logic Display~
6 860 85 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 QB
-6 -32 8 -24
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89727e-315 5.42414e-315
0
14 Logic Display~
6 800 86 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 QD
-10 -32 4 -24
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89727e-315 5.41896e-315
0
14 Logic Display~
6 830 86 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 QC
-5 -33 9 -25
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89727e-315 5.41378e-315
0
9 Inverter~
13 812 172 0 2 22
0 4 25
0
0 0 608 90
6 74LS04
-15 31 27 39
3 U5A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7168 0 0
2
5.89727e-315 5.4086e-315
0
9 Inverter~
13 842 173 0 2 22
0 17 32
0
0 0 608 90
6 74LS04
-11 38 31 46
3 U5B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3171 0 0
2
5.89727e-315 5.40342e-315
0
9 Inverter~
13 872 173 0 2 22
0 18 31
0
0 0 608 90
6 74LS04
3 32 45 40
3 U5C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4139 0 0
2
5.89727e-315 5.39824e-315
0
10 3-In NAND~
219 550 110 0 4 22
0 25 17 18 48
0
0 0 608 0
6 74LS10
2 -33 44 -25
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 5 0
1 U
6435 0 0
2
5.89727e-315 5.39306e-315
0
10 3-In NAND~
219 550 156 0 4 22
0 25 28 33 47
0
0 0 608 0
6 74LS10
10 -34 52 -26
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
5283 0 0
2
5.89727e-315 5.38788e-315
0
10 3-In NAND~
219 550 256 0 4 22
0 32 18 28 45
0
0 0 608 0
6 74LS10
6 -36 48 -28
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 5 0
1 U
6874 0 0
2
5.89727e-315 5.37752e-315
0
10 3-In NAND~
219 550 205 0 4 22
0 25 32 28 46
0
0 0 608 0
6 74LS10
5 -34 47 -26
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
5305 0 0
2
5.89727e-315 5.36716e-315
0
10 2-In NAND~
219 555 307 0 3 22
0 4 28 44
0
0 0 608 0
4 7400
6 -36 34 -28
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
34 0 0
2
5.89727e-315 5.3568e-315
0
10 2-In NAND~
219 555 355 0 3 22
0 4 17 43
0
0 0 608 0
4 7400
11 -37 39 -29
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
969 0 0
2
5.89727e-315 5.34643e-315
0
10 3-In NAND~
219 553 410 0 4 22
0 17 18 28 42
0
0 0 608 0
6 74LS10
-2 -35 40 -27
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
8402 0 0
2
5.89727e-315 5.32571e-315
0
10 3-In NAND~
219 555 457 0 4 22
0 17 31 27 41
0
0 0 608 0
6 74LS10
5 -35 47 -27
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 6 0
1 U
3751 0 0
2
5.89727e-315 5.30499e-315
0
10 4-In NAND~
219 654 170 0 5 22
0 48 47 46 45 30
0
0 0 608 0
6 74LS20
-27 -39 15 -31
4 U11A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
4292 0 0
2
5.89727e-315 5.26354e-315
0
10 4-In NAND~
219 653 382 0 5 22
0 44 43 42 41 29
0
0 0 608 0
6 74LS20
-21 -28 21 -20
4 U11B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
6118 0 0
2
5.89727e-315 0
0
7 74LS154
95 1054 168 0 22 45
0 2 2 16 4 17 18 64 65 66
67 68 69 70 71 6 7 8 72 9
10 73 74
0
0 0 4832 0
7 74LS154
-27 -98 22 -90
2 U1
-7 -88 7 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.89727e-315 0
0
91
1 0 3 0 0 4096 0 23 0 0 20 2
1166 82
1166 96
1 0 4 0 0 4096 0 9 0 0 17 2
925 149
925 276
3 2 5 0 0 12416 0 21 9 0 0 4
951 176
951 163
943 163
943 149
15 1 6 0 0 8320 0 54 16 0 0 4
1092 177
1112 177
1112 144
1143 144
16 1 7 0 0 4224 0 54 15 0 0 4
1092 186
1122 186
1122 180
1144 180
17 1 8 0 0 4224 0 54 13 0 0 4
1092 195
1124 195
1124 213
1144 213
19 1 9 0 0 8320 0 54 14 0 0 4
1092 213
1111 213
1111 248
1145 248
20 1 10 0 0 8320 0 54 12 0 0 4
1092 222
1100 222
1100 284
1145 284
2 1 11 0 0 4224 0 12 11 0 0 3
1181 284
1425 284
1425 80
2 1 12 0 0 4224 0 14 10 0 0 3
1181 248
1373 248
1373 83
2 1 13 0 0 4224 0 13 17 0 0 3
1180 213
1331 213
1331 83
2 1 14 0 0 4224 0 15 18 0 0 3
1180 180
1288 180
1288 85
2 1 15 0 0 4224 0 16 19 0 0 3
1179 144
1244 144
1244 82
0 2 2 0 0 8192 0 0 54 15 0 3
997 148
997 159
1016 159
1 1 2 0 0 4096 0 20 54 0 0 3
997 120
997 150
1016 150
0 3 16 0 0 8320 0 0 54 91 0 5
800 253
800 292
989 292
989 186
1022 186
0 4 4 0 0 8192 0 0 54 90 0 5
829 244
829 276
1000 276
1000 195
1022 195
0 5 17 0 0 8192 0 0 54 22 0 4
960 259
1009 259
1009 204
1022 204
0 6 18 0 0 4096 0 0 54 21 0 4
942 241
1018 241
1018 213
1022 213
3 1 3 0 0 8320 0 9 22 0 0 6
934 103
934 57
1115 57
1115 96
1204 96
1204 82
0 1 18 0 0 0 0 0 21 88 0 4
889 226
889 241
942 241
942 222
0 2 17 0 0 8192 0 0 21 89 0 4
859 235
859 259
960 259
960 222
1 6 19 0 0 20608 0 36 26 0 0 8
706 181
683 181
683 193
638 193
638 283
390 283
390 438
278 438
4 3 20 0 0 4224 0 27 26 0 0 2
186 456
230 456
2 1 21 0 0 8320 0 26 1 0 0 4
230 438
219 438
219 399
187 399
1 4 22 0 0 4224 0 24 26 0 0 2
254 508
254 486
1 1 23 0 0 4224 0 26 25 0 0 2
254 411
254 397
6 1 24 0 0 4224 0 36 28 0 0 3
700 253
659 253
659 242
0 9 25 0 0 4096 0 0 36 73 0 3
774 148
774 199
770 199
7 0 2 0 0 0 0 36 0 0 31 3
770 181
786 181
786 190
8 0 2 0 0 0 0 36 0 0 32 3
770 190
786 190
786 208
10 0 2 0 0 8320 0 36 0 0 33 4
770 208
786 208
786 287
737 287
4 1 2 0 0 0 0 36 29 0 0 5
706 226
670 226
670 287
739 287
739 303
5 3 26 0 0 8320 0 36 30 0 0 4
706 235
694 235
694 512
580 512
0 2 27 0 0 4096 0 0 30 39 0 3
493 466
493 521
534 521
0 1 28 0 0 4096 0 0 30 42 0 3
503 419
503 503
534 503
5 3 29 0 0 8320 0 53 36 0 0 4
680 382
683 382
683 208
706 208
5 2 30 0 0 8320 0 52 36 0 0 4
681 170
693 170
693 199
706 199
0 3 27 0 0 8320 0 0 51 55 0 3
333 338
333 466
531 466
2 2 31 0 0 20608 0 43 51 0 0 7
875 155
875 129
751 129
751 50
444 50
444 457
531 457
0 1 17 0 0 0 0 0 51 44 0 3
492 401
492 448
531 448
0 3 28 0 0 4096 0 0 50 47 0 3
503 314
503 419
529 419
0 2 18 0 0 4096 0 0 50 50 0 3
471 256
471 410
529 410
0 1 17 0 0 0 0 0 50 45 0 3
492 364
492 401
529 401
0 2 17 0 0 12288 0 0 49 72 0 5
502 108
502 148
492 148
492 364
531 364
0 1 4 0 0 0 0 0 49 48 0 3
458 298
458 346
531 346
0 2 28 0 0 0 0 0 48 49 0 3
503 265
503 316
531 316
0 1 4 0 0 0 0 0 48 85 0 3
458 128
458 298
531 298
0 3 28 0 0 0 0 0 46 52 0 3
503 214
503 265
526 265
0 2 18 0 0 4096 0 0 46 87 0 3
471 20
471 256
526 256
0 1 32 0 0 8192 0 0 46 53 0 3
481 205
481 247
526 247
0 3 28 0 0 0 0 0 47 56 0 3
503 156
503 214
526 214
2 2 32 0 0 16512 0 42 47 0 0 7
845 155
845 139
739 139
739 61
481 61
481 205
526 205
2 3 33 0 0 12416 0 31 45 0 0 5
333 287
333 267
433 267
433 165
526 165
13 1 27 0 0 0 0 33 31 0 0 5
290 285
309 285
309 338
333 338
333 323
13 2 28 0 0 4224 0 32 45 0 0 4
291 175
416 175
416 156
526 156
0 1 25 0 0 0 0 0 47 58 0 3
512 147
512 196
526 196
0 1 25 0 0 0 0 0 45 73 0 3
512 101
512 147
526 147
0 5 17 0 0 0 0 0 33 86 0 5
355 139
355 211
219 211
219 303
226 303
0 6 18 0 0 0 0 0 33 87 0 5
345 148
345 203
210 203
210 312
226 312
11 1 2 0 0 0 0 33 35 0 0 5
296 267
310 267
310 216
331 216
331 225
9 1 2 0 0 0 0 32 34 0 0 5
297 121
313 121
313 70
334 70
334 79
0 2 34 0 0 4224 0 0 33 66 0 3
190 148
190 276
226 276
1 1 35 0 0 4224 0 6 33 0 0 4
115 325
180 325
180 267
226 267
3 1 36 0 0 4224 0 32 2 0 0 4
227 139
143 139
143 99
119 99
4 1 34 0 0 0 0 32 3 0 0 4
227 148
134 148
134 136
115 136
1 5 37 0 0 12416 0 5 32 0 0 5
114 176
134 176
134 159
227 159
227 157
1 6 38 0 0 12416 0 4 32 0 0 4
117 212
142 212
142 166
227 166
1 7 39 0 0 12416 0 8 32 0 0 4
115 249
148 249
148 175
227 175
1 8 40 0 0 8320 0 7 32 0 0 4
116 288
154 288
154 184
227 184
0 3 18 0 0 0 0 0 44 87 0 3
490 20
490 119
526 119
0 2 17 0 0 0 0 0 44 86 0 3
502 28
502 110
526 110
2 1 25 0 0 16512 0 41 44 0 0 7
815 154
815 148
729 148
729 70
512 70
512 101
526 101
0 1 18 0 0 0 0 0 43 88 0 3
890 198
875 198
875 191
0 1 17 0 0 0 0 0 42 89 0 3
860 199
845 199
845 191
0 1 4 0 0 0 0 0 41 90 0 3
830 198
815 198
815 190
4 4 41 0 0 8320 0 51 53 0 0 4
582 457
602 457
602 396
629 396
3 4 42 0 0 4224 0 53 50 0 0 4
629 387
593 387
593 410
580 410
3 2 43 0 0 12416 0 49 53 0 0 4
582 355
593 355
593 378
629 378
3 1 44 0 0 8320 0 48 53 0 0 4
582 307
601 307
601 369
629 369
4 4 45 0 0 8320 0 46 52 0 0 4
577 256
601 256
601 184
630 184
4 3 46 0 0 12416 0 47 52 0 0 4
577 205
593 205
593 175
630 175
4 2 47 0 0 12416 0 45 52 0 0 4
577 156
592 156
592 166
630 166
4 1 48 0 0 8320 0 44 52 0 0 4
577 110
601 110
601 157
630 157
0 10 4 0 0 12416 0 0 32 90 0 7
830 120
814 120
814 35
458 35
458 129
291 129
291 130
0 11 17 0 0 12416 0 0 32 89 0 6
860 119
843 119
843 28
434 28
434 139
291 139
0 12 18 0 0 12416 0 0 32 88 0 6
890 120
875 120
875 20
415 20
415 148
291 148
11 1 18 0 0 0 0 36 37 0 0 3
770 226
890 226
890 103
12 1 17 0 0 0 0 36 38 0 0 3
770 235
860 235
860 103
13 1 4 0 0 0 0 36 40 0 0 3
770 244
830 244
830 104
14 1 16 0 0 0 0 36 39 0 0 3
770 253
800 253
800 104
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
