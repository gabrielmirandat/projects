CircuitMaker Text
5.6
Probes: 5
R3_2
AC Analysis
0 344 255 65280
R3_2
DC Sweep
0 344 255 65280
R3_2
Operating Point
0 344 255 65280
R3_2
Fourier Analysis
0 344 255 65280
V2_1
Transient Analysis
0 249 254 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 200 5 100 10
176 79 1364 455
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
93 C:\Users\Marina\Documents\4� semestre\Sistemas digitais 1\Laborat�rio\CircuitMakerfim\BOM.DAT
0 7
2 2 0.386943 0.500000
344 175 1532 418
9961490 0
0
6 Title:
5 Name:
0
0
0
6
5 SAVE-
218 344 255 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
5130 0 0
2
42269 0
0
7 Ground~
168 322 336 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
42269 1
0
11 Signal Gen~
195 208 280 0 19 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1084227584
20
1 1000 0 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -5/5V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 5 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
42269 2
0
9 Resistor~
219 322 285 0 3 5
0 2 3 -1
0
0 0 880 90
7 1000000
-9 0 40 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
3421 0 0
2
5.89724e-315 0
0
9 Resistor~
219 388 283 0 3 5
0 2 3 -1
0
0 0 880 90
6 100.13
-6 0 36 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8157 0 0
2
42269 3
0
9 Resistor~
219 279 255 0 2 5
0 4 3
0
0 0 880 0
2 50
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
5572 0 0
2
42269 4
0
6
0 1 2 0 0 4096 0 0 2 2 0 2
322 308
322 330
0 1 2 0 0 4096 0 0 5 5 0 3
321 308
388 308
388 301
0 2 3 0 0 4224 0 0 5 4 0 3
322 255
388 255
388 265
2 2 3 0 0 0 0 6 4 0 0 3
297 255
322 255
322 267
2 1 2 0 0 12416 0 3 4 0 0 5
239 285
242 285
242 308
322 308
322 303
1 1 4 0 0 8320 0 3 6 0 0 4
239 275
242 275
242 255
261 255
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
