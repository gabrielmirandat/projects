CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1550 0 3 120 10
176 79 1364 707
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
93 C:\Users\Marina\Documents\4� semestre\Sistemas digitais 1\Laborat�rio\CircuitMakerfim\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
58
13 Logic Switch~
5 782 147 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6869 0 0
2
41929.7 0
0
13 Logic Switch~
5 781 52 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
952 0 0
2
41929.7 1
0
10 2-In NAND~
219 1682 214 0 3 22
0 33 3 4
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
522 0 0
2
5.89681e-315 0
0
10 2-In NAND~
219 1687 343 0 3 22
0 7 32 10
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
733 0 0
2
5.89681e-315 0
0
9 Inverter~
13 1740 389 0 2 22
0 11 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U18A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
6533 0 0
2
5.89681e-315 0
0
9 Inverter~
13 145 226 0 2 22
0 17 16
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
8922 0 0
2
5.89681e-315 0
0
10 StopLight~
181 2027 374 0 12 13
0 18 4 5 0 0 0 0 0 0
2 2 2
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM2
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
3391 0 0
2
41929.7 2
0
10 StopLight~
181 1974 238 0 12 13
0 19 10 12 0 0 0 0 0 0
2 2 2
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM1
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
342 0 0
2
41929.7 3
0
5 7425~
219 304 276 0 6 22
0 23 24 22 25 20 21
0
0 0 608 0
4 7425
-14 -24 14 -16
3 U9A
-3 19 18 27
0
15 DVCC=14;DGND=7;
69 %D [%14bi %7bi %1i %2i %3i %4i %5i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 5 4 2 1 3 6 5 4 2
1 3 6 9 10 12 13 11 8 0
0 6 0
65 0 0 0 2 1 7 0
1 U
4297 0 0
2
41929.7 4
0
7 Ground~
168 403 449 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8118 0 0
2
41929.7 5
0
2 +V
167 429 345 0 1 3
0 26
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V16
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3254 0 0
2
41929.7 6
0
7 74LS160
124 524 382 0 14 29
0 26 26 21 16 2 2 2 2 26
69 28 27 14 15
0
0 0 4832 0
7 74LS160
-24 -51 25 -43
2 U1
-8 -52 6 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3562 0 0
2
41929.7 7
0
9 2-In AND~
219 110 226 0 3 22
0 19 18 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
4351 0 0
2
41929.7 8
0
2 +V
167 174 64 0 1 3
0 29
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V15
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6645 0 0
2
41929.7 9
0
7 Ground~
168 183 202 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9648 0 0
2
41929.7 10
0
7 74LS160
124 215 144 0 14 29
0 29 29 30 16 2 70 71 72 29
73 23 24 22 25
0
0 0 4832 0
7 74LS160
-24 -51 25 -43
3 U17
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
358 0 0
2
41929.7 11
0
2 +V
167 1797 389 0 1 3
0 31
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V14
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5822 0 0
2
41929.7 12
0
10 8-In NAND~
219 1842 441 0 9 19
0 9 11 7 31 31 31 32 8 18
0
0 0 608 0
6 74LS30
-21 -24 21 -16
3 U16
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
3905 0 0
2
41929.7 13
0
2 +V
167 1636 182 0 1 3
0 13
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V13
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
853 0 0
2
41929.7 14
0
10 8-In NAND~
219 1676 290 0 9 19
0 33 3 6 8 13 13 13 9 19
0
0 0 608 0
6 74LS30
-21 -24 21 -16
3 U15
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
8452 0 0
2
41929.7 15
0
9 Inverter~
13 1276 364 0 2 22
0 74 75
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U14F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 6 9 0
1 U
7616 0 0
2
41929.7 16
0
9 Inverter~
13 1302 324 0 2 22
0 76 77
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U14E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 5 9 0
1 U
3445 0 0
2
41929.7 17
0
9 Inverter~
13 1359 382 0 2 22
0 78 79
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U14D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 4 9 0
1 U
6281 0 0
2
41929.7 18
0
9 Inverter~
13 1790 530 0 2 22
0 6 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
8532 0 0
2
41929.7 19
0
7 Ground~
168 1491 337 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7947 0 0
2
41929.7 20
0
2 +V
167 1462 287 0 1 3
0 34
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V12
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3620 0 0
2
41929.7 21
0
7 74LS138
19 1535 286 0 14 29
0 35 36 37 34 2 2 33 3 6
8 32 7 11 9
0
0 0 5088 0
7 74LS138
-25 -61 24 -53
3 U13
-11 -71 10 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5855 0 0
2
41929.7 22
0
9 Inverter~
13 1592 106 0 2 22
0 39 38
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 U6D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
7464 0 0
2
41929.7 23
0
2 +V
167 1462 61 0 1 3
0 40
0
0 0 54240 0
3 10V
-11 -22 10 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6374 0 0
2
41929.7 24
0
7 Ground~
168 1123 152 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3957 0 0
2
41929.7 25
0
14 Logic Display~
6 1507 126 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3702 0 0
2
41929.7 26
0
14 Logic Display~
6 1482 115 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9398 0 0
2
41929.7 27
0
14 Logic Display~
6 1467 108 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6929 0 0
2
41929.7 28
0
9 3-In AND~
219 1538 134 0 4 22
0 35 36 37 39
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 3 0
1 U
6608 0 0
2
41929.7 29
0
9 2-In AND~
219 842 139 0 3 22
0 47 48 45
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
7927 0 0
2
41929.7 30
0
9 2-In AND~
219 837 62 0 3 22
0 49 47 46
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3378 0 0
2
41929.7 31
0
8 2-In OR~
219 919 148 0 3 22
0 45 44 42
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
7964 0 0
2
41929.7 32
0
8 2-In OR~
219 914 67 0 3 22
0 46 44 43
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
5711 0 0
2
41929.7 33
0
2 +V
167 998 105 0 1 3
0 50
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3105 0 0
2
41929.7 34
0
7 74LS151
20 1064 192 0 14 29
0 50 50 43 50 50 50 42 50 2
35 36 37 41 80
0
0 0 4832 0
7 74LS151
-24 -60 25 -52
3 U11
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3951 0 0
2
41929.7 35
0
7 74LS161
96 1425 106 0 14 29
0 41 41 30 81 82 83 84 40 38
85 86 35 36 37
0
0 0 4832 0
8 74LS161A
-28 -60 28 -52
3 U10
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3274 0 0
2
41929.7 36
0
14 Logic Display~
6 662 503 0 1 2
10 44
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9252 0 0
2
5.89681e-315 0
0
9 2-In AND~
219 593 520 0 3 22
0 15 14 44
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4860 0 0
2
5.89681e-315 5.26354e-315
0
2 +V
167 502 13 0 1 3
0 51
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3282 0 0
2
5.89681e-315 5.30499e-315
0
5 7474~
219 538 66 0 6 22
0 51 51 59 16 87 47
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
9535 0 0
2
5.89681e-315 5.32571e-315
0
14 Logic Display~
6 629 13 0 1 2
10 47
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5822 0 0
2
5.89681e-315 5.34643e-315
0
9 Inverter~
13 328 57 0 2 22
0 22 60
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3155 0 0
2
5.89681e-315 5.3568e-315
0
9 3-In AND~
219 395 48 0 4 22
0 24 60 25 59
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
9153 0 0
2
5.89681e-315 5.36716e-315
0
4 4511
219 666 427 0 14 29
0 28 27 14 15 2 61 61 52 53
54 55 56 57 58
0
0 0 4832 0
4 4511
-14 -60 14 -52
2 U5
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
9839 0 0
2
41929.7 37
0
2 +V
167 608 460 0 1 3
0 61
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3277 0 0
2
41929.7 38
0
7 Ground~
168 535 463 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
372 0 0
2
41929.7 39
0
9 CC 7-Seg~
183 614 173 0 16 19
10 58 57 56 55 54 53 52 2 2
2 2 2 2 2 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
782 0 0
2
41929.7 40
0
7 Ground~
168 578 121 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9330 0 0
2
41929.7 41
0
9 CC 7-Seg~
183 508 173 0 16 19
10 62 63 68 67 66 65 64 2 2
2 2 2 2 2 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
797 0 0
2
41929.7 42
0
7 Ground~
168 227 225 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7896 0 0
2
41929.7 43
0
2 +V
167 300 222 0 1 3
0 20
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3527 0 0
2
41929.7 44
0
4 4511
219 358 189 0 20 29
0 23 24 22 25 2 20 20 64 65
66 67 68 63 62 0 0 0 0 0
5
0
0 0 4832 0
4 4511
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7535 0 0
2
41929.7 45
0
7 Pulser~
4 74 153 0 10 12
0 88 89 30 90 0 0 10 10 11
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7444 0 0
2
41929.7 46
0
154
0 2 3 0 0 4096 0 0 3 68 0 3
1613 268
1613 223
1658 223
3 0 4 0 0 0 0 3 0 0 62 2
1709 214
1709 214
2 3 5 0 0 4224 0 24 7 0 0 4
1811 530
1991 530
1991 388
2011 388
1 0 6 0 0 0 0 24 0 0 5 2
1775 530
1775 530
0 0 6 0 0 4224 0 0 0 69 0 3
1580 277
1580 530
1779 530
0 3 7 0 0 8320 0 0 18 9 0 3
1647 334
1647 428
1818 428
0 8 8 0 0 8320 0 0 18 70 0 3
1607 286
1607 473
1818 473
0 1 9 0 0 8320 0 0 18 71 0 3
1638 322
1638 410
1818 410
12 1 7 0 0 0 0 27 4 0 0 4
1573 304
1625 304
1625 334
1663 334
3 0 10 0 0 0 0 4 0 0 64 2
1714 343
1714 343
0 2 11 0 0 8320 0 0 18 13 0 3
1701 389
1701 419
1818 419
2 3 12 0 0 4224 0 5 8 0 0 4
1761 389
1926 389
1926 252
1958 252
13 1 11 0 0 0 0 27 5 0 0 4
1573 313
1616 313
1616 389
1725 389
0 7 13 0 0 8192 0 0 20 15 0 3
1636 304
1636 313
1652 313
0 6 13 0 0 0 0 0 20 16 0 3
1636 295
1636 304
1652 304
1 5 13 0 0 4224 0 19 20 0 0 3
1636 191
1636 295
1652 295
13 2 14 0 0 4224 0 12 43 0 0 3
556 409
556 529
569 529
0 1 15 0 0 4224 0 0 43 44 0 3
562 418
562 511
569 511
2 4 16 0 0 4096 0 6 16 0 0 3
166 226
166 144
177 144
4 2 16 0 0 4096 0 12 6 0 0 3
486 382
166 382
166 226
1 3 17 0 0 4224 0 6 13 0 0 2
130 226
131 226
4 0 16 0 0 4224 0 45 0 0 19 4
538 78
152 78
152 160
166 160
0 2 18 0 0 8320 0 0 13 57 0 5
1903 441
1903 649
67 649
67 235
86 235
0 1 19 0 0 4096 0 0 13 25 0 4
623 619
42 619
42 217
86 217
0 0 19 0 0 4096 0 0 0 26 0 2
1301 619
619 619
0 0 19 0 0 16512 0 0 0 66 0 5
1893 290
1893 180
2104 180
2104 619
1292 619
0 2 4 0 0 8320 0 0 7 62 0 3
1841 214
1841 374
2011 374
0 1 18 0 0 0 0 0 7 57 0 3
1954 441
1954 360
2011 360
0 5 20 0 0 8192 0 0 9 149 0 3
310 238
309 238
309 255
6 0 21 0 0 0 0 9 0 0 36 2
343 276
343 276
3 0 22 0 0 4096 0 9 0 0 39 2
287 281
288 281
8 0 2 0 0 4096 0 12 0 0 35 2
492 418
403 418
7 0 2 0 0 0 0 12 0 0 35 2
492 409
403 409
6 0 2 0 0 0 0 12 0 0 35 2
492 400
403 400
1 5 2 0 0 0 0 10 12 0 0 3
403 443
403 391
492 391
0 3 21 0 0 12416 0 0 12 0 0 4
335 276
344 276
344 373
492 373
0 1 23 0 0 4224 0 0 9 137 0 3
254 153
254 263
287 263
0 2 24 0 0 4096 0 0 9 136 0 3
270 162
270 272
287 272
0 0 22 0 0 4096 0 0 0 135 0 3
288 171
288 281
293 281
0 4 25 0 0 4224 0 0 9 134 0 3
279 180
279 290
287 290
9 0 26 0 0 8320 0 12 0 0 43 4
562 355
562 319
461 319
461 354
2 1 26 0 0 0 0 12 11 0 0 3
492 364
429 364
429 354
1 1 26 0 0 0 0 12 11 0 0 3
492 355
492 354
429 354
4 14 15 0 0 0 0 49 12 0 0 2
634 418
556 418
3 13 14 0 0 0 0 49 12 0 0 2
634 409
556 409
2 12 27 0 0 4224 0 49 12 0 0 2
634 400
556 400
1 11 28 0 0 4224 0 49 12 0 0 2
634 391
556 391
0 9 29 0 0 4224 0 0 16 50 0 4
174 98
262 98
262 117
253 117
0 2 29 0 0 0 0 0 16 50 0 3
174 117
174 126
183 126
1 1 29 0 0 0 0 14 16 0 0 3
174 73
174 117
183 117
5 1 2 0 0 0 0 16 15 0 0 2
183 153
183 196
3 3 30 0 0 4096 0 58 16 0 0 4
98 144
159 144
159 135
183 135
14 0 25 0 0 0 0 16 0 0 134 2
247 180
247 180
13 0 22 0 0 0 0 16 0 0 135 2
247 171
247 171
12 0 24 0 0 0 0 16 0 0 136 2
247 162
247 162
11 0 23 0 0 0 0 16 0 0 137 2
247 153
247 153
9 0 18 0 0 0 0 18 0 0 0 2
1869 441
1959 441
0 6 31 0 0 8192 0 0 18 59 0 3
1797 446
1797 455
1818 455
0 5 31 0 0 0 0 0 18 60 0 3
1797 437
1797 446
1818 446
1 4 31 0 0 4224 0 17 18 0 0 3
1797 398
1797 437
1818 437
0 7 32 0 0 8320 0 0 18 65 0 3
1657 352
1657 464
1818 464
0 0 4 0 0 0 0 0 0 0 0 2
1705 214
1857 214
0 1 33 0 0 8320 0 0 3 67 0 3
1577 259
1577 205
1658 205
0 2 10 0 0 4224 0 0 8 0 0 4
1710 343
1949 343
1949 238
1958 238
11 2 32 0 0 0 0 27 4 0 0 4
1573 295
1586 295
1586 352
1663 352
9 1 19 0 0 0 0 20 8 0 0 4
1703 290
1935 290
1935 224
1958 224
7 1 33 0 0 0 0 27 20 0 0 2
1573 259
1652 259
8 2 3 0 0 4224 0 27 20 0 0 2
1573 268
1652 268
9 3 6 0 0 0 0 27 20 0 0 2
1573 277
1652 277
10 4 8 0 0 0 0 27 20 0 0 2
1573 286
1652 286
14 8 9 0 0 0 0 27 20 0 0 2
1573 322
1652 322
6 0 2 0 0 0 0 27 0 0 73 2
1497 322
1491 322
5 1 2 0 0 0 0 27 25 0 0 3
1497 313
1491 313
1491 331
1 4 34 0 0 8320 0 26 27 0 0 3
1462 296
1462 304
1503 304
0 1 35 0 0 4096 0 0 27 90 0 3
1459 174
1459 259
1503 259
0 2 36 0 0 4096 0 0 27 89 0 3
1444 183
1444 268
1503 268
0 3 37 0 0 4096 0 0 27 88 0 3
1429 192
1429 277
1503 277
2 9 38 0 0 8320 0 28 41 0 0 3
1595 88
1595 79
1463 79
4 1 39 0 0 4224 0 34 28 0 0 3
1559 134
1595 134
1595 124
1 8 40 0 0 4224 0 29 41 0 0 2
1462 70
1463 70
9 1 2 0 0 0 0 40 30 0 0 3
1102 165
1102 146
1123 146
1 0 37 0 0 0 0 31 0 0 85 2
1507 144
1507 143
1 0 36 0 0 0 0 32 0 0 86 2
1482 133
1482 133
1 0 35 0 0 0 0 33 0 0 90 2
1467 126
1467 124
0 3 37 0 0 0 0 0 34 88 0 3
1472 145
1472 143
1514 143
2 0 36 0 0 0 0 34 0 0 89 3
1514 134
1514 133
1482 133
0 1 35 0 0 0 0 0 34 90 0 3
1499 124
1499 125
1514 125
14 12 37 0 0 12416 0 41 40 0 0 4
1457 142
1472 142
1472 192
1096 192
13 11 36 0 0 12416 0 41 40 0 0 4
1457 133
1482 133
1482 183
1096 183
12 10 35 0 0 12416 0 41 40 0 0 4
1457 124
1499 124
1499 174
1096 174
2 0 41 0 0 4096 0 41 0 0 92 2
1393 79
1369 79
13 1 41 0 0 4224 0 40 41 0 0 4
1096 219
1369 219
1369 70
1393 70
3 7 42 0 0 8320 0 37 40 0 0 3
952 148
952 219
1032 219
3 3 43 0 0 8320 0 38 40 0 0 4
947 67
973 67
973 183
1032 183
0 2 44 0 0 4096 0 0 37 110 0 2
895 157
906 157
3 1 45 0 0 4224 0 35 37 0 0 2
863 139
906 139
3 1 46 0 0 4224 0 36 38 0 0 3
858 62
901 62
901 58
0 1 47 0 0 4096 0 0 35 123 0 3
792 71
792 130
818 130
1 2 48 0 0 8320 0 1 35 0 0 3
794 147
794 148
818 148
1 1 49 0 0 8320 0 2 36 0 0 3
793 52
793 53
813 53
6 0 50 0 0 4096 0 40 0 0 105 2
1032 210
998 210
5 0 50 0 0 0 0 40 0 0 105 2
1032 201
998 201
4 0 50 0 0 0 0 40 0 0 105 2
1032 192
998 192
2 0 50 0 0 0 0 40 0 0 105 2
1032 174
998 174
0 8 50 0 0 4224 0 0 40 106 0 3
998 165
998 228
1032 228
1 1 50 0 0 0 0 39 40 0 0 3
998 114
998 165
1032 165
0 3 30 0 0 8320 0 0 41 52 0 3
128 144
128 88
1393 88
0 1 19 0 0 0 0 0 13 0 0 3
80 204
80 217
86 217
1 0 44 0 0 0 0 42 0 0 110 2
662 521
662 520
3 2 44 0 0 8320 0 43 38 0 0 4
614 520
895 520
895 76
901 76
2 1 51 0 0 4224 0 45 45 0 0 3
514 30
514 3
538 3
8 7 52 0 0 8320 0 49 52 0 0 5
698 445
742 445
742 295
629 295
629 209
9 6 53 0 0 12416 0 49 52 0 0 5
698 436
787 436
787 281
623 281
623 209
10 5 54 0 0 12416 0 49 52 0 0 5
698 427
827 427
827 234
617 234
617 209
11 4 55 0 0 8320 0 49 52 0 0 5
698 418
802 418
802 223
611 223
611 209
12 3 56 0 0 8320 0 49 52 0 0 5
698 409
729 409
729 263
605 263
605 209
13 2 57 0 0 12416 0 49 52 0 0 5
698 400
758 400
758 251
599 251
599 209
14 1 58 0 0 8320 0 49 52 0 0 5
698 391
705 391
705 231
593 231
593 209
0 8 2 0 0 8320 0 0 52 121 0 5
614 105
642 105
642 213
635 213
635 209
8 0 2 0 0 0 0 54 0 0 140 3
529 209
537 209
537 105
0 9 2 0 0 0 0 0 52 140 0 3
578 105
614 105
614 131
1 0 47 0 0 0 0 46 0 0 123 2
629 31
629 30
6 2 47 0 0 12416 0 45 36 0 0 4
562 30
665 30
665 71
813 71
1 2 51 0 0 0 0 44 45 0 0 5
502 22
502 30
515 30
515 30
514 30
4 3 59 0 0 4224 0 48 45 0 0 2
416 48
514 48
2 2 60 0 0 8320 0 47 48 0 0 3
349 57
349 48
371 48
0 1 22 0 0 4224 0 0 47 135 0 2
313 171
313 57
0 3 25 0 0 0 0 0 48 134 0 5
320 180
320 122
367 122
367 57
371 57
0 1 24 0 0 4224 0 0 48 136 0 3
303 162
303 39
371 39
0 7 61 0 0 8192 0 0 49 133 0 3
618 439
618 445
628 445
5 1 2 0 0 0 0 49 51 0 0 5
628 427
576 427
576 440
535 440
535 457
7 7 61 0 0 0 0 49 49 0 0 4
628 445
628 440
628 440
628 445
6 1 61 0 0 8320 0 49 50 0 0 5
628 436
618 436
618 477
608 477
608 469
4 0 25 0 0 0 0 57 0 0 0 2
326 180
244 180
3 0 22 0 0 0 0 57 0 0 0 2
326 171
244 171
2 0 24 0 0 0 0 57 0 0 0 2
326 162
244 162
0 1 23 0 0 0 0 0 57 0 0 2
244 153
326 153
14 1 62 0 0 4224 0 57 54 0 0 5
390 153
477 153
477 227
487 227
487 209
13 2 63 0 0 8320 0 57 54 0 0 5
390 162
463 162
463 255
493 255
493 209
9 1 2 0 0 0 0 54 53 0 0 4
508 131
508 105
578 105
578 115
7 0 64 0 0 0 0 54 0 0 150 2
523 209
523 209
6 0 65 0 0 0 0 54 0 0 151 2
517 209
517 209
5 0 66 0 0 0 0 54 0 0 152 2
511 209
511 209
4 0 67 0 0 0 0 54 0 0 153 2
505 209
505 209
3 0 68 0 0 0 0 54 0 0 154 2
499 209
499 209
0 7 20 0 0 0 0 0 57 149 0 3
310 201
310 207
320 207
5 1 2 0 0 0 0 57 55 0 0 5
320 189
268 189
268 202
227 202
227 219
7 7 20 0 0 0 0 57 57 0 0 4
320 207
320 202
320 202
320 207
6 1 20 0 0 8320 0 57 56 0 0 5
320 198
310 198
310 239
300 239
300 231
8 0 64 0 0 12416 0 57 0 0 0 5
390 207
396 207
396 333
523 333
523 206
9 0 65 0 0 8320 0 57 0 0 0 5
390 198
401 198
401 324
517 324
517 206
10 0 66 0 0 8320 0 57 0 0 0 5
390 189
408 189
408 312
511 312
511 206
11 0 67 0 0 8320 0 57 0 0 0 5
390 180
417 180
417 295
505 295
505 206
12 0 68 0 0 8320 0 57 0 0 0 5
390 171
431 171
431 267
499 267
499 206
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2017 318 2114 339
2025 325 2105 340
10 SEMAFOROEW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1956 183 2061 204
1964 190 2052 205
11 SEMAFORO NS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1798 193 1881 214
1807 200 1871 215
8 EWYELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1901 420 1958 441
1909 427 1949 442
5 EWRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1752 326 1833 347
1760 332 1824 347
8 NSYELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1804 506 1877 527
1812 513 1868 528
7 EWGREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1698 347 1773 368
1707 353 1763 368
7 NSGREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1714 271 1771 292
1722 277 1762 292
5 NSRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
768 157 827 178
777 163 817 178
5 ewcar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
762 7 819 28
770 14 810 29
5 nscar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
81 247 138 268
89 253 129 268
5 ewred
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
94 181 151 202
102 187 142 202
5 nsred
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
456 118 537 139
464 125 528 140
8 unidades
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
649 127 722 148
657 133 713 148
7 dezenas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
671 13 744 34
679 20 735 35
7 TMSHORT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
738 462 805 483
747 469 795 484
6 TMLONG
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
