CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
23 C:\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 1532 489
9469970 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 97 279 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6857 0 0
2
42187 0
0
13 Logic Switch~
5 95 228 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
428 0 0
2
42187 0
0
13 Logic Switch~
5 94 174 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6131 0 0
2
42187 0
0
9 Inverter~
13 239 352 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
9516 0 0
2
42187 0
0
10 2-In NAND~
219 642 262 0 3 22
0 2 12 3
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4529 0 0
2
42187 0
0
10 2-In NAND~
219 638 179 0 3 22
0 13 3 2
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4226 0 0
2
42187 0
0
10 2-In NAND~
219 501 265 0 3 22
0 4 9 12
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3561 0 0
2
42187 0
0
10 2-In NAND~
219 500 177 0 3 22
0 8 4 13
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
368 0 0
2
42187 0
0
10 2-In NAND~
219 348 265 0 3 22
0 8 10 9
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
386 0 0
2
42187 0
0
10 2-In NAND~
219 350 177 0 3 22
0 11 9 8
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6544 0 0
2
42187 0
0
10 3-In NAND~
219 236 270 0 4 22
0 5 6 2 10
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
8869 0 0
2
42187 0
0
10 3-In NAND~
219 237 174 0 4 22
0 3 7 5 11
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
3573 0 0
2
42187 0
0
14 Logic Display~
6 896 137 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7945 0 0
2
42187 0
0
14 Logic Display~
6 840 137 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6306 0 0
2
42187 0
0
21
3 0 2 0 0 8320 0 11 0 0 21 4
212 279
212 390
828 390
828 179
1 0 3 0 0 12416 0 12 0 0 20 5
213 165
172 165
172 92
757 92
757 262
2 0 4 0 0 4240 0 4 0 0 13 4
260 352
452 352
452 219
477 219
0 1 5 0 0 4224 0 0 4 5 0 3
149 228
149 352
224 352
1 0 5 0 0 0 0 2 0 0 6 2
107 228
212 228
3 1 5 0 0 0 0 12 11 0 0 3
213 183
212 183
212 261
1 2 6 0 0 4224 0 1 11 0 0 4
109 279
193 279
193 270
212 270
1 2 7 0 0 4224 0 3 12 0 0 2
106 174
213 174
0 1 8 0 0 8192 0 0 9 17 0 5
386 177
386 223
297 223
297 256
324 256
2 0 9 0 0 12416 0 10 0 0 16 5
326 186
295 186
295 210
396 210
396 265
4 2 10 0 0 4224 0 11 9 0 0 4
263 270
316 270
316 274
324 274
4 1 11 0 0 4224 0 12 10 0 0 4
264 174
318 174
318 168
326 168
2 1 4 0 0 0 0 8 7 0 0 3
476 186
477 186
477 256
1 0 2 0 0 0 0 5 0 0 21 5
618 253
590 253
590 225
684 225
684 179
2 0 3 0 0 0 0 6 0 0 20 5
614 188
589 188
589 215
718 215
718 262
3 2 9 0 0 0 0 9 7 0 0 4
375 265
469 265
469 274
477 274
3 1 8 0 0 4224 0 10 8 0 0 4
377 177
468 177
468 168
476 168
3 2 12 0 0 4224 0 7 5 0 0 4
528 265
610 265
610 271
618 271
3 1 13 0 0 4224 0 8 6 0 0 4
527 177
606 177
606 170
614 170
3 1 3 0 0 0 0 5 13 0 0 3
669 262
896 262
896 155
3 1 2 0 0 0 0 6 14 0 0 3
665 179
840 179
840 155
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
879 86 916 110
889 94 905 110
2 QB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
824 86 853 110
834 94 842 110
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
49 215 78 239
59 223 67 239
1 T
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
49 263 78 287
59 271 67 287
1 K
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
49 160 78 184
59 168 67 184
1 J
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
