CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
43037874 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 30 241 0 1 11
0 40
0
0 0 22368 0
2 0V
-7 -18 7 -10
1 Z
-3 -28 4 -20
8 AUXILIAR
-27 -36 29 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
6770 0 0
2
42248.9 0
0
13 Logic Switch~
5 41 871 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
3 V10
-10 -28 11 -20
1 D
-3 -36 4 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3305 0 0
2
42248.9 1
0
13 Logic Switch~
5 41 822 0 1 11
0 16
0
0 0 21856 0
2 0V
-7 -18 7 -10
2 V9
-7 -28 7 -20
1 C
-3 -36 4 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5643 0 0
2
42248.9 2
0
13 Logic Switch~
5 41 776 0 1 11
0 17
0
0 0 21856 0
2 0V
-7 -18 7 -10
2 V8
-7 -28 7 -20
1 B
-3 -36 4 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8224 0 0
2
42248.9 3
0
13 Logic Switch~
5 42 728 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
2 V7
-7 -28 7 -20
1 A
-3 -36 4 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6752 0 0
2
42248.9 4
0
13 Logic Switch~
5 41 521 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
2 V1
-7 -28 7 -20
5 RESET
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7272 0 0
2
42248.9 5
0
13 Logic Switch~
5 92 103 0 1 11
0 38
0
0 0 21856 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
12 CLOCK MANUAL
-41 -36 43 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7364 0 0
2
42248.9 6
0
14 Logic Display~
6 585 753 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3161 0 0
2
42248.9 7
0
9 Inverter~
13 270 701 0 2 22
0 6 5
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U6E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
8131 0 0
2
42248.9 8
0
9 Inverter~
13 268 737 0 2 22
0 8 7
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
6931 0 0
2
42248.9 9
0
9 Inverter~
13 267 772 0 2 22
0 10 9
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
3294 0 0
2
42248.9 10
0
9 Inverter~
13 266 808 0 2 22
0 11 3
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
7630 0 0
2
42248.9 11
0
7 Ground~
168 438 674 0 1 3
0 2
0
0 0 53344 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
358 0 0
2
42248.9 12
0
7 Ground~
168 97 675 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5880 0 0
2
42248.9 13
0
7 74LS151
20 376 752 0 14 29
0 3 7 41 9 3 5 42 9 2
14 13 12 4 43
0
0 0 4832 0
6 74F151
-21 -60 21 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
8118 0 0
2
42248.9 14
0
7 74LS154
95 150 746 0 22 45
0 2 2 18 17 16 15 44 45 46
47 48 49 50 51 52 53 6 54 8
55 10 11
0
0 0 4832 0
6 74F154
-21 -87 21 -79
2 U7
-7 -88 7 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
3174 0 0
2
42248.9 15
0
9 Inverter~
13 114 314 0 2 22
0 4 19
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
5740 0 0
2
5.89721e-315 0
0
9 3-In AND~
219 243 484 0 4 22
0 4 13 25 21
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 5 0
1 U
4612 0 0
2
5.89721e-315 5.26354e-315
0
9 3-In AND~
219 936 296 0 4 22
0 14 13 12 31
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
3929 0 0
2
5.89721e-315 5.30499e-315
0
8 2-In OR~
219 388 192 0 3 22
0 19 23 29
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6505 0 0
2
5.89721e-315 5.32571e-315
0
8 2-In OR~
219 387 143 0 3 22
0 28 24 30
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8290 0 0
2
5.89721e-315 5.34643e-315
0
9 2-In AND~
219 244 418 0 3 22
0 4 14 22
0
0 0 2656 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3585 0 0
2
5.89721e-315 5.3568e-315
0
9 2-In AND~
219 244 353 0 3 22
0 13 27 23
0
0 0 2656 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3540 0 0
2
5.89721e-315 5.36716e-315
0
9 2-In AND~
219 243 284 0 3 22
0 4 26 24
0
0 0 2656 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3422 0 0
2
5.89721e-315 5.37752e-315
0
9 2-In AND~
219 243 227 0 3 22
0 4 12 28
0
0 0 2656 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4464 0 0
2
5.89721e-315 5.38788e-315
0
14 Logic Display~
6 692 409 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3396 0 0
2
5.89721e-315 5.39306e-315
0
14 Logic Display~
6 662 412 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
766 0 0
2
5.89721e-315 5.39824e-315
0
2 +V
167 600 401 0 1 3
0 33
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5236 0 0
2
5.89721e-315 5.40342e-315
0
6 74112~
219 600 484 0 7 32
0 33 21 20 19 32 27 12
0
0 0 4704 0
5 74112
4 -60 39 -52
5 FFJK3
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
5714 0 0
2
5.89721e-315 5.4086e-315
0
6 74112~
219 602 332 0 7 32
0 34 22 20 19 32 26 13
0
0 0 4704 0
5 74112
4 -60 39 -52
5 FFJK2
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 6 0
1 U
3851 0 0
2
42248.9 16
0
6 74112~
219 603 179 0 7 32
0 35 30 20 29 32 25 14
0
0 0 4704 0
5 74112
4 -60 39 -52
5 FFJK1
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 6 0
1 U
3233 0 0
2
42248.9 17
0
14 Logic Display~
6 684 241 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Q0b
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4890 0 0
2
42248.9 18
0
14 Logic Display~
6 687 98 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Q1b
-11 -20 10 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8536 0 0
2
42248.9 19
0
14 Logic Display~
6 654 242 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5339 0 0
2
42248.9 20
0
14 Logic Display~
6 663 98 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3766 0 0
2
42248.9 21
0
2 +V
167 602 252 0 1 3
0 34
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9987 0 0
2
42248.9 22
0
2 +V
167 602 95 0 1 3
0 35
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9314 0 0
2
42248.9 23
0
14 Logic Display~
6 972 136 0 1 2
10 31
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 S
20 -26 27 -18
6 TRANCA
-21 -41 21 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3502 0 0
2
42248.9 24
0
14 Logic Display~
6 359 52 0 1 2
10 20
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
5 CLOCK
-18 -41 17 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4694 0 0
2
42248.9 25
0
7 Pulser~
4 82 157 0 10 12
0 37 56 36 57 0 0 2 2 2
8
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7703 0 0
2
42248.9 26
0
2 +V
167 228 186 0 1 3
0 39
0
0 0 54240 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
365 0 0
2
42248.9 27
0
2 +V
167 227 43 0 1 3
0 37
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
37 0 0
2
42248.9 28
0
5 7474~
219 227 139 0 6 22
0 37 38 36 39 58 20
0
0 0 864 0
4 7474
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
8938 0 0
2
42248.9 29
0
68
5 0 3 0 0 4096 0 15 0 0 10 2
344 761
333 761
13 1 4 0 0 4096 0 15 8 0 0 3
408 779
585 779
585 771
6 2 5 0 0 8320 0 15 9 0 0 4
344 770
321 770
321 701
291 701
17 1 6 0 0 8320 0 16 9 0 0 4
188 773
216 773
216 701
255 701
2 2 7 0 0 4224 0 10 15 0 0 4
289 737
327 737
327 734
344 734
19 1 8 0 0 8320 0 16 10 0 0 4
188 791
227 791
227 737
253 737
4 0 9 0 0 8192 0 15 0 0 8 3
344 752
327 752
327 788
2 8 9 0 0 8320 0 11 15 0 0 3
288 772
288 788
344 788
21 1 10 0 0 4224 0 16 11 0 0 4
188 809
236 809
236 772
252 772
2 1 3 0 0 8320 0 12 15 0 0 4
287 808
333 808
333 725
344 725
22 1 11 0 0 4224 0 16 12 0 0 4
188 818
243 818
243 808
251 808
0 12 12 0 0 4096 0 0 15 42 0 3
486 538
486 752
408 752
0 11 13 0 0 4096 0 0 15 36 0 3
472 567
472 743
408 743
0 10 14 0 0 4096 0 0 15 32 0 3
459 596
459 734
408 734
9 1 2 0 0 8192 0 15 13 0 0 3
414 725
438 725
438 682
1 0 2 0 0 0 0 16 0 0 17 2
112 728
97 728
1 2 2 0 0 4224 0 14 16 0 0 3
97 683
97 737
112 737
1 6 15 0 0 8320 0 2 16 0 0 4
53 871
88 871
88 791
118 791
1 5 16 0 0 8320 0 3 16 0 0 4
53 822
83 822
83 782
118 782
1 4 17 0 0 12416 0 4 16 0 0 4
53 776
82 776
82 773
118 773
1 3 18 0 0 8320 0 5 16 0 0 4
54 728
83 728
83 764
118 764
0 4 19 0 0 8192 0 0 29 25 0 3
303 314
303 466
576 466
0 3 20 0 0 4096 0 0 29 55 0 3
544 305
544 457
570 457
4 2 21 0 0 12416 0 18 29 0 0 4
264 484
343 484
343 448
576 448
4 0 19 0 0 4224 0 30 0 0 28 2
578 314
303 314
2 3 22 0 0 4224 0 30 22 0 0 4
578 296
329 296
329 418
265 418
3 2 23 0 0 8320 0 23 20 0 0 4
265 353
315 353
315 201
375 201
2 1 19 0 0 0 0 17 20 0 0 4
135 314
303 314
303 183
375 183
2 3 24 0 0 8320 0 21 24 0 0 4
374 152
291 152
291 284
264 284
1 0 4 0 0 0 0 17 0 0 38 2
99 314
74 314
0 3 25 0 0 12416 0 0 18 58 0 6
686 161
843 161
843 609
125 609
125 493
219 493
0 2 14 0 0 8320 0 0 22 46 0 5
802 143
802 596
139 596
139 427
220 427
0 1 13 0 0 0 0 0 23 36 0 3
170 485
170 344
220 344
1 0 4 0 0 0 0 22 0 0 38 2
220 409
74 409
0 2 26 0 0 12416 0 0 24 57 0 6
684 314
762 314
762 582
155 582
155 293
219 293
0 2 13 0 0 8320 0 0 18 37 0 5
724 296
724 567
170 567
170 484
219 484
0 2 13 0 0 0 0 0 19 60 0 2
653 296
912 296
0 1 4 0 0 4096 0 0 18 40 0 3
74 275
74 475
219 475
2 0 27 0 0 12416 0 23 0 0 49 5
220 362
185 362
185 552
692 552
692 465
1 0 4 0 0 0 0 24 0 0 41 2
219 275
74 275
1 0 4 0 0 20608 0 25 0 0 2 7
219 218
74 218
74 275
16 275
16 631
524 631
524 779
2 0 12 0 0 12416 0 25 0 0 47 5
219 236
199 236
199 538
662 538
662 448
3 1 28 0 0 12416 0 25 21 0 0 4
264 227
280 227
280 134
374 134
4 3 29 0 0 4224 0 31 20 0 0 4
579 161
448 161
448 192
421 192
2 3 30 0 0 4224 0 31 21 0 0 2
579 143
420 143
0 1 14 0 0 0 0 0 19 61 0 4
663 143
892 143
892 287
912 287
0 3 12 0 0 0 0 0 19 50 0 4
662 448
893 448
893 305
912 305
4 1 31 0 0 8320 0 19 38 0 0 3
957 296
972 296
972 154
1 6 27 0 0 0 0 26 29 0 0 3
692 427
692 466
630 466
7 1 12 0 0 0 0 29 27 0 0 3
624 448
662 448
662 430
5 0 32 0 0 8192 0 29 0 0 56 3
600 496
600 521
503 521
1 1 33 0 0 4224 0 28 29 0 0 2
600 410
600 421
5 0 32 0 0 8192 0 30 0 0 56 3
602 344
602 355
503 355
1 1 34 0 0 4224 0 36 30 0 0 2
602 261
602 269
0 3 20 0 0 0 0 0 30 59 0 3
544 200
544 305
572 305
5 1 32 0 0 16512 0 31 6 0 0 5
603 191
603 210
503 210
503 521
53 521
6 1 26 0 0 0 0 30 32 0 0 3
632 314
684 314
684 259
6 1 25 0 0 0 0 31 33 0 0 3
633 161
687 161
687 116
0 3 20 0 0 4224 0 0 31 63 0 6
359 103
544 103
544 200
544 200
544 152
573 152
7 1 13 0 0 0 0 30 34 0 0 3
626 296
654 296
654 260
7 1 14 0 0 0 0 31 35 0 0 3
627 143
663 143
663 116
1 1 35 0 0 4224 0 37 31 0 0 4
602 104
602 126
603 126
603 116
6 1 20 0 0 0 0 43 39 0 0 3
251 103
359 103
359 70
3 3 36 0 0 12416 0 40 43 0 0 4
106 148
151 148
151 121
203 121
0 1 37 0 0 4224 0 0 40 68 0 4
227 59
28 59
28 148
58 148
1 2 38 0 0 4224 0 7 43 0 0 2
104 103
203 103
4 1 39 0 0 4224 0 43 41 0 0 3
227 151
227 171
228 171
1 1 37 0 0 0 0 42 43 0 0 2
227 52
227 76
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
