CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 210 10
238 79 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
34 C:\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
406 175 519 272
42991634 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 232 184 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 Enable
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
336 0 0
2
42152.9 0
0
13 Logic Switch~
5 36 27 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
618 0 0
2
42152.9 0
0
13 Logic Switch~
5 36 295 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5663 0 0
2
42152.9 1
0
13 Logic Switch~
5 34 260 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
367 0 0
2
42152.9 2
0
13 Logic Switch~
5 33 224 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8112 0 0
2
42152.9 3
0
13 Logic Switch~
5 34 188 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4359 0 0
2
42152.9 4
0
13 Logic Switch~
5 34 149 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
855 0 0
2
42152.9 5
0
13 Logic Switch~
5 35 108 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3572 0 0
2
42152.9 6
0
13 Logic Switch~
5 34 62 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7676 0 0
2
42152.9 7
0
14 Logic Display~
6 327 121 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 GotNoth
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3645 0 0
2
42152.9 8
0
14 Logic Display~
6 476 122 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3275 0 0
2
42152.9 9
0
14 Logic Display~
6 454 122 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
979 0 0
2
42152.9 10
0
14 Logic Display~
6 433 123 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3481 0 0
2
42152.9 11
0
9 Inverter~
13 390 300 0 2 22
0 9 4
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
6542 0 0
2
42152.9 12
0
9 Inverter~
13 390 273 0 2 22
0 10 5
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3361 0 0
2
42152.9 13
0
9 Inverter~
13 390 248 0 2 22
0 11 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9647 0 0
2
42152.9 14
0
9 Inverter~
13 389 223 0 2 22
0 12 7
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8891 0 0
2
42152.9 15
0
9 Inverter~
13 387 196 0 2 22
0 13 8
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8581 0 0
2
42152.9 16
0
14 Logic Display~
6 270 119 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 GotSome
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7669 0 0
2
42152.9 17
0
5 74148
219 310 232 0 14 29
0 2 3 16 17 18 19 15 14 20
9 10 11 12 13
0
0 0 4848 0
5 74148
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 3 2 1 13 12 11 10
15 9 7 6 14 5 4 3 2 1
13 12 11 10 15 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
367 0 0
2
42152.9 19
0
28
1 1 2 0 0 4224 0 1 20 0 0 4
244 184
264 184
264 196
272 196
1 7 3 0 0 4096 0 2 0 0 28 4
48 27
66 27
66 43
84 43
1 2 4 0 0 20608 0 10 14 0 0 7
327 139
327 154
416 154
416 90
495 90
495 300
411 300
2 1 5 0 0 8320 0 15 11 0 0 3
411 273
476 273
476 140
1 2 6 0 0 4224 0 12 16 0 0 3
454 140
454 248
411 248
2 1 7 0 0 8320 0 17 13 0 0 3
410 223
433 223
433 141
2 1 8 0 0 12416 0 18 19 0 0 5
408 196
420 196
420 163
270 163
270 137
10 1 9 0 0 8320 0 20 14 0 0 4
348 277
356 277
356 300
375 300
11 1 10 0 0 8320 0 20 15 0 0 4
348 241
362 241
362 273
375 273
12 1 11 0 0 4224 0 20 16 0 0 4
348 232
371 232
371 248
375 248
1 13 12 0 0 4224 0 17 20 0 0 2
374 223
348 223
14 1 13 0 0 4224 0 20 18 0 0 2
348 196
372 196
1 1 14 0 0 8192 0 0 4 28 0 4
84 289
64 289
64 260
46 260
1 2 15 0 0 12288 0 5 0 0 28 4
45 224
57 224
57 202
84 202
3 6 16 0 0 4224 0 20 0 0 28 2
272 223
84 223
7 2 15 0 0 4224 0 20 0 0 28 2
272 259
84 259
4 5 17 0 0 4224 0 20 0 0 28 2
272 232
84 232
5 4 18 0 0 4224 0 20 0 0 28 2
272 241
84 241
6 3 19 0 0 4224 0 20 0 0 28 2
272 250
84 250
8 1 14 0 0 4224 0 20 0 0 28 2
272 268
84 268
9 0 20 0 0 4224 0 20 0 0 28 2
272 277
84 277
2 7 3 0 0 4224 0 20 0 0 28 2
272 214
84 214
1 6 16 0 0 0 0 9 0 0 28 2
46 62
84 62
1 5 17 0 0 0 0 8 0 0 28 2
47 108
84 108
1 4 18 0 0 0 0 7 0 0 28 2
46 149
84 149
1 3 19 0 0 0 0 6 0 0 28 2
46 188
84 188
1 0 20 0 0 0 0 3 0 0 28 2
48 295
84 295
-46 0 1 0 0 4256 0 0 0 0 0 2
84 29
84 324
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
