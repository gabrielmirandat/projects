CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9469970 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 42 272 0 1 11
0 13
0
0 0 22368 0
2 0V
-6 -16 8 -8
1 M
-3 -26 4 -18
5 MOEDA
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3710 0 0
2
42243.6 0
0
13 Logic Switch~
5 244 521 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
2 V1
-7 -28 7 -20
5 RESET
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3931 0 0
2
42243.6 1
0
13 Logic Switch~
5 92 103 0 1 11
0 20
0
0 0 21856 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
12 CLOCK MANUAL
-41 -36 43 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3696 0 0
2
42243.6 2
0
9 2-In AND~
219 832 360 0 3 22
0 5 4 2
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3143 0 0
2
42243.6 3
0
9 2-In AND~
219 831 191 0 3 22
0 5 6 3
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3245 0 0
2
42243.6 4
0
9 Inverter~
13 60 357 0 2 22
0 13 10
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U4A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
980 0 0
2
42243.6 5
0
8 2-In OR~
219 221 390 0 3 22
0 10 4 9
0
0 0 2656 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4848 0 0
2
42243.6 6
0
8 2-In OR~
219 222 300 0 3 22
0 13 6 12
0
0 0 608 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6220 0 0
2
42243.6 7
0
9 2-In AND~
219 440 325 0 3 22
0 8 9 7
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5603 0 0
2
42243.6 8
0
14 Logic Display~
6 684 386 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Q0b
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3873 0 0
2
42243.6 9
0
14 Logic Display~
6 683 141 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Q1b
-11 -20 10 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3521 0 0
2
42243.6 10
0
9 2-In AND~
219 440 260 0 3 22
0 8 12 11
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
393 0 0
2
42243.6 11
0
14 Logic Display~
6 652 388 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4578 0 0
2
42243.6 12
0
14 Logic Display~
6 651 143 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3283 0 0
2
42243.6 13
0
2 +V
167 602 348 0 1 3
0 15
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3919 0 0
2
42243.6 14
0
2 +V
167 602 102 0 1 3
0 16
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8669 0 0
2
42243.6 15
0
14 Logic Display~
6 971 283 0 1 2
10 2
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 E
20 -26 27 -18
4 ERRO
-14 -41 14 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8151 0 0
2
42243.6 16
0
14 Logic Display~
6 972 136 0 1 2
10 3
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 R
20 -26 27 -18
7 RETORNO
-24 -41 25 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
524 0 0
2
42243.6 17
0
14 Logic Display~
6 359 52 0 1 2
10 17
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
5 CLOCK
-18 -41 17 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4926 0 0
2
42243.6 18
0
7 Pulser~
4 82 157 0 10 12
0 19 22 18 23 0 0 2 2 10
8
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5600 0 0
2
42243.6 19
0
2 +V
167 228 215 0 1 3
0 21
0
0 0 54240 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8789 0 0
2
42243.6 20
0
2 +V
167 227 31 0 1 3
0 19
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9673 0 0
2
42243.6 21
0
5 7474~
219 602 474 0 6 22
0 15 7 17 14 4 6
0
0 0 4704 0
4 7474
7 -60 35 -52
2 D0
25 -61 39 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 1 2 0
1 U
647 0 0
2
42243.6 22
0
5 7474~
219 602 227 0 6 22
0 16 11 17 14 8 5
0
0 0 4704 0
4 7474
7 -60 35 -52
2 D1
25 -61 39 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 0 2 2 1 0
1 U
3847 0 0
2
42243.6 23
0
5 7474~
219 227 139 0 6 22
0 19 20 18 21 24 17
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3449 0 0
2
42243.6 24
0
33
3 1 2 0 0 4224 0 4 17 0 0 3
853 360
971 360
971 301
3 1 3 0 0 4224 0 5 18 0 0 3
852 191
972 191
972 154
0 2 4 0 0 4096 0 0 4 10 0 4
684 457
775 457
775 369
808 369
0 1 5 0 0 4224 0 0 4 6 0 3
652 191
652 351
808 351
0 2 6 0 0 8192 0 0 5 12 0 4
652 438
714 438
714 200
807 200
0 1 5 0 0 0 0 0 5 21 0 4
650 191
749 191
749 182
807 182
3 2 7 0 0 8320 0 9 23 0 0 4
461 325
500 325
500 438
578 438
0 1 8 0 0 4096 0 0 9 14 0 3
398 250
398 316
416 316
3 2 9 0 0 4224 0 7 9 0 0 4
254 390
399 390
399 334
416 334
0 2 4 0 0 8320 0 0 7 18 0 5
684 456
684 586
95 586
95 399
208 399
2 1 10 0 0 8320 0 6 7 0 0 3
63 375
63 381
208 381
0 2 6 0 0 8320 0 0 8 20 0 5
652 438
652 555
140 555
140 309
209 309
3 2 11 0 0 4224 0 12 24 0 0 4
461 260
530 260
530 191
578 191
0 1 8 0 0 8320 0 0 12 19 0 7
683 209
683 254
505 254
505 196
398 196
398 251
416 251
3 2 12 0 0 12416 0 8 12 0 0 4
255 300
324 300
324 269
416 269
0 1 13 0 0 4224 0 0 8 17 0 2
63 291
209 291
1 1 13 0 0 0 0 1 6 0 0 3
54 272
63 272
63 339
5 1 4 0 0 0 0 23 10 0 0 3
632 456
684 456
684 404
5 1 8 0 0 0 0 24 11 0 0 3
632 209
683 209
683 159
6 1 6 0 0 0 0 23 13 0 0 3
626 438
652 438
652 406
6 1 5 0 0 0 0 24 14 0 0 3
626 191
651 191
651 161
4 0 14 0 0 12288 0 24 0 0 23 4
602 239
602 293
523 293
523 521
1 4 14 0 0 4224 0 2 23 0 0 3
256 521
602 521
602 486
1 1 15 0 0 4224 0 15 23 0 0 2
602 357
602 411
1 1 16 0 0 4224 0 16 24 0 0 2
602 111
602 164
0 3 17 0 0 4224 0 0 23 27 0 3
564 209
564 456
578 456
0 3 17 0 0 0 0 0 24 28 0 4
359 103
564 103
564 209
578 209
6 1 17 0 0 0 0 25 19 0 0 3
251 103
359 103
359 70
3 3 18 0 0 12416 0 20 25 0 0 4
106 148
151 148
151 121
203 121
0 1 19 0 0 4224 0 0 20 33 0 4
227 48
28 48
28 148
58 148
1 2 20 0 0 4224 0 3 25 0 0 2
104 103
203 103
4 1 21 0 0 4224 0 25 21 0 0 3
227 151
227 200
228 200
1 1 19 0 0 0 0 22 25 0 0 2
227 40
227 76
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
