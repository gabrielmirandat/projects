CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
328 139 1343 676
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
496 235 609 332
43024530 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 49 182 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9672 0 0
2
5.89725e-315 0
0
2 +V
167 152 20 0 1 3
0 3
0
0 0 54256 0
3 10V
4 -8 25 0
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
42276 0
0
2 +V
167 153 137 0 1 3
0 4
0
0 0 54256 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6369 0 0
2
5.89725e-315 0
0
5 7474~
219 152 99 0 6 22
0 3 6 2 4 19 5
0
0 0 4720 0
4 7474
9 -70 37 -62
3 U6A
14 -61 35 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
9172 0 0
2
5.89725e-315 0
0
7 Pulser~
4 46 128 0 10 12
0 3 20 2 21 0 0 10 10 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7100 0 0
2
5.89725e-315 0
0
9 2-In XOR~
219 802 340 0 3 22
0 7 9 8
0
0 0 112 0
5 74F86
-13 -31 22 -23
3 U5A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3820 0 0
2
42276 0
0
8 2-In OR~
219 500 303 0 3 22
0 12 11 10
0
0 0 112 0
5 74F32
-14 -31 21 -23
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7678 0 0
2
42276 1
0
8 2-In OR~
219 577 353 0 3 22
0 10 16 9
0
0 0 112 0
5 74F32
-12 -30 23 -22
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
961 0 0
2
42276 2
0
8 2-In OR~
219 570 228 0 3 22
0 13 14 7
0
0 0 112 0
5 74F32
-11 -35 24 -27
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3178 0 0
2
42276 3
0
9 2-In AND~
219 397 390 0 3 22
0 17 9 11
0
0 0 112 0
5 74F08
-21 -28 14 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3409 0 0
2
42276 4
0
9 2-In AND~
219 398 328 0 3 22
0 5 17 12
0
0 0 112 0
5 74F08
-23 -27 12 -19
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3951 0 0
2
42276 5
0
9 2-In AND~
219 401 266 0 3 22
0 5 7 14
0
0 0 112 0
5 74F08
-23 -25 12 -17
3 U2C
-7 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8885 0 0
2
5.89725e-315 5.26354e-315
0
14 Logic Display~
6 859 158 0 1 2
10 7
0
0 0 53856 0
6 100MEG
-21 -33 21 -25
1 D
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89725e-315 5.30499e-315
0
14 Logic Display~
6 863 308 0 1 2
10 8
0
0 0 53856 0
6 100MEG
-24 -35 18 -27
1 M
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.89725e-315 5.32571e-315
0
9 Inverter~
13 483 480 0 2 22
0 7 17
0
0 0 368 180
5 74F04
-13 -25 22 -17
3 U1B
-5 -30 16 -22
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9442 0 0
2
5.89725e-315 5.34643e-315
0
14 Logic Display~
6 644 287 0 1 2
10 9
0
0 0 53856 0
6 100MEG
-20 -32 22 -24
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89725e-315 5.3568e-315
0
9 2-In AND~
219 403 214 0 3 22
0 7 9 15
0
0 0 112 0
5 74F08
-24 -28 11 -20
3 U2B
-15 -24 6 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9968 0 0
2
5.89725e-315 5.36716e-315
0
14 Logic Display~
6 636 167 0 1 2
10 7
0
0 0 53856 0
6 100MEG
-20 -32 22 -24
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89725e-315 5.37752e-315
0
8 2-In OR~
219 489 184 0 3 22
0 16 15 13
0
0 0 112 0
5 74F32
-13 -29 22 -21
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8464 0 0
2
5.89725e-315 5.38788e-315
0
9 2-In AND~
219 400 157 0 3 22
0 18 9 16
0
0 0 112 0
5 74F08
-22 -31 13 -23
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7168 0 0
2
5.89725e-315 5.39306e-315
0
9 Inverter~
13 143 243 0 2 22
0 5 18
0
0 0 368 0
5 74F04
-17 -27 18 -19
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3171 0 0
2
5.89725e-315 5.39824e-315
0
31
3 3 2 0 0 12416 0 5 4 0 0 4
70 119
86 119
86 81
128 81
1 0 3 0 0 12416 0 5 0 0 3 4
22 119
10 119
10 31
152 31
1 1 3 0 0 0 0 2 4 0 0 2
152 29
152 36
1 4 4 0 0 8320 0 3 4 0 0 3
153 122
152 122
152 111
1 0 5 0 0 4096 0 21 0 0 24 2
128 243
120 243
1 2 6 0 0 8320 0 1 4 0 0 4
61 182
103 182
103 63
128 63
0 1 7 0 0 4096 0 0 13 28 0 3
738 228
859 228
859 176
3 1 8 0 0 4224 0 6 14 0 0 3
835 340
863 340
863 326
0 2 9 0 0 4096 0 0 6 27 0 4
644 355
772 355
772 349
786 349
1 0 7 0 0 0 0 6 0 0 28 2
786 331
738 331
3 1 10 0 0 8320 0 7 8 0 0 4
533 303
547 303
547 344
564 344
2 3 11 0 0 8320 0 7 10 0 0 4
487 312
480 312
480 390
418 390
3 1 12 0 0 4224 0 11 7 0 0 4
419 328
462 328
462 294
487 294
3 1 13 0 0 8320 0 19 9 0 0 4
522 184
536 184
536 219
557 219
3 2 14 0 0 12416 0 12 9 0 0 4
422 266
462 266
462 237
557 237
3 2 15 0 0 4224 0 17 19 0 0 4
424 214
461 214
461 193
476 193
0 2 16 0 0 4224 0 0 8 18 0 3
446 175
446 362
564 362
3 1 16 0 0 0 0 20 19 0 0 4
421 157
446 157
446 175
476 175
2 0 9 0 0 4096 0 10 0 0 27 2
373 399
216 399
1 0 17 0 0 4096 0 10 0 0 22 2
373 381
255 381
0 1 5 0 0 8192 0 0 11 24 0 3
120 257
120 319
374 319
2 2 17 0 0 4224 0 15 11 0 0 4
468 480
255 480
255 337
374 337
2 0 7 0 0 4096 0 12 0 0 26 2
377 275
235 275
6 1 5 0 0 20608 0 4 12 0 0 6
176 63
194 63
194 135
120 135
120 257
377 257
2 0 9 0 0 4096 0 17 0 0 27 2
379 223
216 223
0 1 7 0 0 12416 0 0 17 28 0 5
537 480
537 510
235 510
235 205
379 205
0 2 9 0 0 8320 0 0 20 30 0 5
644 353
644 529
216 529
216 166
376 166
0 1 7 0 0 0 0 0 15 29 0 4
635 228
738 228
738 480
504 480
3 1 7 0 0 0 0 9 18 0 0 3
603 228
636 228
636 185
3 1 9 0 0 0 0 8 16 0 0 3
610 353
644 353
644 305
2 1 18 0 0 12416 0 21 20 0 0 4
164 243
186 243
186 148
376 148
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
