CircuitMaker Text
5.6
Probes: 8
C_2
AC Analysis
1 392 87 65535
C_2
DC Sweep
1 392 87 65535
C_2
Fourier Analysis
1 392 87 65535
V2_1
AC Analysis
0 198 87 65280
V2_1
DC Sweep
0 198 87 65280
V2_1
Operating Point
0 198 87 65280
V2_1
Fourier Analysis
0 198 87 65280
L_2
Transient Analysis
0 398 87 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 1 1
20 Package,Description,
93 C:\Users\Marina\Documents\4� semestre\Sistemas digitais 1\Laborat�rio\CircuitMakerfim\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 1532 489
1083703314 0
0
6 Title:
5 Name:
0
0
0
7
5 SAVE-
218 392 87 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
7361 0 0
2
5.89731e-315 0
0
5 SAVE-
218 198 87 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4747 0 0
2
5.89731e-315 5.26354e-315
0
9 Inductor~
219 352 87 0 2 5
0 4 3
0
0 0 848 0
7 1.05 mH
-24 -17 25 -9
1 L
-4 -27 3 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89731e-315 5.30499e-315
0
7 Ground~
168 297 216 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
5.89731e-315 5.32571e-315
0
10 Capacitor~
219 426 139 0 2 5
0 2 3
0
0 0 848 90
8 0.927 nF
-1 3 55 11
1 C
18 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9998 0 0
2
5.89731e-315 5.34643e-315
0
11 Signal Gen~
195 116 142 0 64 64
0 5 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182400512 -1073741824 1073741824
0 814313567 814313567 939725423 948114031 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 62
20
0 16000 -2 2 0 1e-09 1e-09 3.125e-05 6.25e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -2/2V
-17 -30 18 -22
2 V2
-7 -40 7 -32
0
0
46 %D %1 %2 DC 0 PULSE(-2 2 0 1n 1n 31.25u 62.5u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
5.89731e-315 5.3568e-315
0
9 Resistor~
219 243 87 0 2 5
0 5 4
0
0 0 880 0
7 0.532 k
-26 -14 23 -6
1 R
-4 -24 3 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
4597 0 0
2
5.89731e-315 5.36716e-315
0
5
2 2 3 0 0 4224 0 3 5 0 0 3
370 87
426 87
426 130
0 1 2 0 0 4096 0 0 4 4 0 2
297 188
297 210
2 1 4 0 0 4224 0 7 3 0 0 2
261 87
334 87
2 1 2 0 0 12416 0 6 5 0 0 5
147 147
175 147
175 188
426 188
426 148
1 1 5 0 0 8320 0 6 7 0 0 4
147 137
175 137
175 87
225 87
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 4e-05 4e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
