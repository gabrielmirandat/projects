CircuitMaker Text
5.6
Probes: 6
v2#branch
Operating Point
0 235 272 65280
r1[i]
Operating Point
1 296 254 65535
c1[i]
Operating Point
2 323 286 16776960
V2_1
Transient Analysis
0 244 259 65280
R1_2
Transient Analysis
1 305 255 65535
GND
Transient Analysis
2 306 310 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 190 5 100 10
341 118 1356 655
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 1 1
20 Package,Description,
93 C:\Users\Marina\Documents\4� semestre\Sistemas digitais 1\Laborat�rio\CircuitMakerfim\BOM.DAT
0 7
2 4 0.500000 0.500000
509 214 622 311
9961490 0
0
6 Title:
5 Name:
0
0
0
7
5 SAVE-
218 301 308 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 C
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
8402 0 0
2
5.89727e-315 0
0
5 SAVE-
218 306 255 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3751 0 0
2
5.89727e-315 0
0
5 SAVE-
218 249 255 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4292 0 0
2
5.89727e-315 0
0
10 Capacitor~
219 322 282 0 2 5
0 2 3
0
0 0 832 90
5 0.1uF
10 3 45 11
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6118 0 0
2
5.89727e-315 0
0
7 Ground~
168 285 335 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
34 0 0
2
42294.6 0
0
11 Signal Gen~
195 208 280 0 24 64
0 4 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1144753160 -1082130432 1065462268
0 814313567 814313567 976715828 984528911
20
0 750.188 -1 1.013 0 1e-09 1e-09 0.0007 0.001333 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
9 -1/1.013V
-31 -30 32 -22
2 V2
-7 -40 7 -32
0
0
49 %D %1 %2 DC 0 PULSE(-1 1.013 0 1n 1n 700u 1.333m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6357 0 0
2
42294.6 1
0
9 Resistor~
219 279 255 0 2 5
0 4 3
0
0 0 864 0
4 1050
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
319 0 0
2
42294.6 2
0
4
0 1 2 0 0 4096 0 0 5 3 0 2
285 308
285 329
2 2 3 0 0 4224 0 7 4 0 0 3
297 255
322 255
322 273
2 1 2 0 0 12416 0 6 4 0 0 5
239 285
242 285
242 308
322 308
322 291
1 1 4 0 0 8320 0 6 7 0 0 4
239 275
242 275
242 255
261 255
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
