CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 79 1364 384
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
23 C:\CircuitMaker\BOM.DAT
0 7
5 2 0.500000 0.500000
176 393 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 64 170 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
42192 0
0
13 Logic Switch~
5 59 85 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
42192 1
0
5 SCOPE
12 103 219 0 1 11
0 4
0
0 0 57584 0
1 T
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3124 0 0
2
42192 2
0
5 SCOPE
12 94 47 0 1 11
0 3
0
0 0 57584 0
1 J
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3421 0 0
2
5.89713e-315 0
0
5 SCOPE
12 134 46 0 1 11
0 2
0
0 0 57584 0
1 K
-4 -4 3 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8157 0 0
2
5.89713e-315 0
0
5 SCOPE
12 215 152 0 1 11
0 7
0
0 0 57584 0
1 Q
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5572 0 0
2
42192 3
0
7 Pulser~
4 26 125 0 10 12
0 10 11 5 12 0 0 10 10 2
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
42192 4
0
5 SCOPE
12 279 150 0 1 11
0 6
0
0 0 57584 0
2 QB
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7361 0 0
2
42192 5
0
9 Inverter~
13 98 127 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4747 0 0
2
42192 6
0
2 +V
167 148 211 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
42192 7
0
2 +V
167 170 53 0 1 3
0 9
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
42192 8
0
14 Logic Display~
6 299 85 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
42192 9
0
14 Logic Display~
6 250 86 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
42192 10
0
6 74112~
219 169 141 0 7 32
0 9 3 4 2 8 6 7
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
4597 0 0
2
42192 11
0
13
1 0 2 0 0 8320 0 5 0 0 9 5
134 58
121 58
121 165
111 165
111 170
1 0 3 0 0 4096 0 4 0 0 7 2
94 59
94 85
1 0 4 0 0 12416 0 3 0 0 8 5
103 231
103 235
132 235
132 121
126 121
3 1 5 0 0 4224 0 7 9 0 0 4
50 116
75 116
75 127
83 127
1 0 6 0 0 12288 0 8 0 0 10 6
279 162
279 166
301 166
301 128
295 128
295 123
1 0 7 0 0 12416 0 6 0 0 11 4
215 164
215 168
237 168
237 105
1 2 3 0 0 4224 0 2 14 0 0 4
71 85
131 85
131 105
145 105
2 3 4 0 0 0 0 9 14 0 0 4
119 127
126 127
126 114
139 114
1 4 2 0 0 0 0 1 14 0 0 4
76 170
142 170
142 123
145 123
6 1 6 0 0 4224 0 14 12 0 0 3
199 123
299 123
299 103
7 1 7 0 0 0 0 14 13 0 0 5
193 105
238 105
238 112
250 112
250 104
1 5 8 0 0 12416 0 10 14 0 0 4
148 220
148 224
169 224
169 153
1 1 9 0 0 4224 0 11 14 0 0 4
170 62
170 70
169 70
169 78
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
47 91 76 115
57 99 65 115
1 T
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
278 38 315 62
288 46 304 62
2 QB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
236 39 265 63
246 47 254 63
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
22 156 51 180
32 164 40 180
1 K
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
19 70 48 94
29 78 37 94
1 J
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
