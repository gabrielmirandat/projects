* C:\Users\Marina\Desktop\EXP6CBODE.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 27 13:06:57 2015



** Analysis setup **
.ac DEC 101 1K 100K


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EXP6CBODE.net"
.INC "EXP6CBODE.als"


.probe


.END
