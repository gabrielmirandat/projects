CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 740 30 90 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 1 1
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9478322 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 36 194 0 1 11
0 5
0
0 0 21856 0
2 0V
-7 -18 7 -10
2 V7
-7 -28 7 -20
6 ENABLE
-20 -36 22 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89724e-315 0
0
13 Logic Switch~
5 31 305 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 22240 0
2 5V
-7 -18 7 -10
6 UPDOWN
-20 -28 22 -20
7 ENTRADA
-23 -39 26 -31
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89724e-315 5.26354e-315
0
13 Logic Switch~
5 29 523 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -18 7 -10
2 V1
-7 -28 7 -20
5 RESET
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89724e-315 5.30499e-315
0
13 Logic Switch~
5 47 88 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
12 CLOCK MANUAL
-41 -36 43 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89724e-315 5.32571e-315
0
9 2-In AND~
219 109 130 0 3 22
0 7 5 6
0
0 0 2656 0
5 74F08
-18 -36 17 -28
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8157 0 0
2
42269.8 0
0
2 +V
167 871 408 0 1 3
0 8
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
5.89724e-315 5.34643e-315
0
2 +V
167 875 252 0 1 3
0 9
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8901 0 0
2
5.89724e-315 5.3568e-315
0
2 +V
167 876 106 0 1 3
0 10
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89724e-315 5.36716e-315
0
9 Inverter~
13 150 130 0 2 22
0 6 4
0
0 0 608 0
5 74F04
-17 -30 18 -22
3 U8D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
4747 0 0
2
5.89724e-315 5.37752e-315
0
9 Inverter~
13 666 458 0 2 22
0 13 12
0
0 0 608 0
5 74F04
-18 -34 17 -26
3 U8C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
972 0 0
2
5.89724e-315 5.38788e-315
0
9 Inverter~
13 336 322 0 2 22
0 23 22
0
0 0 608 0
5 74F04
-18 -32 17 -24
3 U8B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
3472 0 0
2
42269.8 1
0
9 Inverter~
13 338 261 0 2 22
0 28 27
0
0 0 608 0
5 74F04
-17 -30 18 -22
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
9998 0 0
2
42269.8 2
0
9 2-In XOR~
219 274 492 0 3 22
0 24 25 13
0
0 0 608 0
5 74F86
-18 -24 17 -16
3 U7B
-5 -35 16 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3536 0 0
2
42269.8 3
0
9 2-In XOR~
219 203 460 0 3 22
0 3 16 24
0
0 0 608 0
5 74F86
-18 -35 17 -27
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
4597 0 0
2
42269.8 4
0
9 2-In XOR~
219 210 405 0 3 22
0 3 16 21
0
0 0 608 0
5 74F86
-18 -37 17 -29
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3835 0 0
2
42269.8 5
0
9 2-In XOR~
219 208 339 0 3 22
0 3 16 23
0
0 0 608 0
5 74F86
-18 -35 17 -27
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3670 0 0
2
42269.8 6
0
9 2-In XOR~
219 206 279 0 3 22
0 3 25 28
0
0 0 608 0
5 74F86
-18 -34 17 -26
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5616 0 0
2
42269.8 7
0
9 2-In XOR~
219 205 223 0 3 22
0 3 25 26
0
0 0 608 0
5 74F86
-18 -35 17 -27
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9323 0 0
2
42269.8 8
0
9 3-In AND~
219 1147 296 0 4 22
0 16 15 14 30
0
0 0 608 0
5 74F11
-22 -36 13 -28
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
317 0 0
2
42269.8 9
0
9 2-In AND~
219 471 398 0 3 22
0 21 29 17
0
0 0 2656 0
5 74F08
-20 -37 15 -29
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3108 0 0
2
42269.8 10
0
9 2-In AND~
219 473 331 0 3 22
0 22 29 18
0
0 0 2656 0
5 74F08
-20 -37 15 -29
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4299 0 0
2
42269.8 11
0
9 2-In AND~
219 472 270 0 3 22
0 27 14 19
0
0 0 2656 0
5 74F08
-17 -38 18 -30
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9672 0 0
2
42269.8 12
0
9 2-In AND~
219 471 159 0 3 22
0 26 14 20
0
0 0 2656 0
5 74F08
-18 -36 17 -28
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7876 0 0
2
42269.8 13
0
14 Logic Display~
6 936 413 0 1 2
10 14
0
0 0 53872 0
6 100MEG
0 -34 42 -26
2 Q3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
42269.8 14
0
14 Logic Display~
6 910 411 0 1 2
10 29
0
0 0 53872 0
6 100MEG
-17 -32 25 -24
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
42269.8 15
0
6 74112~
219 871 494 0 7 32
0 8 12 11 13 31 14 29
0
0 0 4704 0
5 74112
-41 -71 -6 -63
5 FFJK3
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
7100 0 0
2
42269.8 16
0
6 74112~
219 876 337 0 7 32
0 9 18 11 17 31 15 25
0
0 0 4704 0
5 74112
-50 -67 -15 -59
5 FFJK2
15 -61 50 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 6 0
1 U
3820 0 0
2
5.89724e-315 5.39306e-315
0
6 74112~
219 876 195 0 7 32
0 10 20 11 19 31 32 16
0
0 0 4704 0
5 74112
4 -60 39 -52
5 FFJK1
-49 -71 -14 -63
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 6 0
1 U
7678 0 0
2
5.89724e-315 5.39824e-315
0
14 Logic Display~
6 981 244 0 1 2
10 15
0
0 0 53872 0
6 100MEG
-54 -30 -12 -22
3 Q0b
-11 -30 10 -22
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89724e-315 5.40342e-315
0
14 Logic Display~
6 1027 102 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -32 45 -24
3 Q1b
26 -20 47 -12
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89724e-315 5.4086e-315
0
14 Logic Display~
6 957 244 0 1 2
10 25
0
0 0 53872 0
6 100MEG
14 -22 56 -14
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89724e-315 5.41378e-315
0
14 Logic Display~
6 1005 102 0 1 2
10 16
0
0 0 53872 0
6 100MEG
-24 -35 18 -27
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.89724e-315 5.41896e-315
0
14 Logic Display~
6 1200 142 0 1 2
10 30
0
0 0 54896 0
6 100MEG
10 -14 52 -6
1 S
20 -26 27 -18
6 ULTIMO
-21 -41 21 -33
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.89724e-315 5.42414e-315
0
14 Logic Display~
6 359 52 0 1 2
10 11
0
0 0 54896 0
6 100MEG
3 -16 45 -8
1 C
-13 -17 -6 -9
5 CLOCK
-9 -29 26 -21
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89724e-315 5.42933e-315
0
7 Pulser~
4 42 130 0 10 12
0 2 35 7 36 0 0 2 2 3
7
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9265 0 0
2
5.89724e-315 5.43192e-315
0
2 +V
167 227 174 0 1 3
0 34
0
0 0 54240 180
3 10V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
5.89724e-315 5.43451e-315
0
2 +V
167 227 46 0 1 3
0 2
0
0 0 54240 0
3 10V
9 -1 30 7
2 V1
14 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9424 0 0
2
5.89724e-315 5.4371e-315
0
5 7474~
219 227 139 0 6 22
0 2 33 4 34 37 11
0
0 0 864 0
4 7474
7 -73 35 -65
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9968 0 0
2
5.89724e-315 5.43969e-315
0
58
1 1 2 0 0 4096 0 38 37 0 0 2
227 76
227 55
1 0 3 0 0 4096 0 17 0 0 41 2
190 270
62 270
1 0 3 0 0 4096 0 16 0 0 5 2
192 330
61 330
1 0 3 0 0 4096 0 15 0 0 5 2
194 396
61 396
0 1 3 0 0 4224 0 0 14 41 0 3
61 305
61 451
187 451
2 3 4 0 0 12416 0 9 38 0 0 4
171 130
177 130
177 121
203 121
2 1 5 0 0 8320 0 5 1 0 0 4
85 139
73 139
73 194
48 194
3 1 6 0 0 4224 0 5 9 0 0 2
130 130
135 130
3 1 7 0 0 4224 0 35 5 0 0 2
66 121
85 121
1 1 8 0 0 4224 0 6 26 0 0 2
871 417
871 431
1 1 9 0 0 4224 0 7 27 0 0 3
875 261
875 274
876 274
1 0 10 0 0 8320 0 8 0 0 54 3
876 115
875 115
875 126
3 0 11 0 0 4096 0 28 0 0 48 2
846 168
807 168
2 2 12 0 0 4224 0 26 10 0 0 2
847 458
687 458
0 1 13 0 0 8192 0 0 10 23 0 3
618 476
618 458
651 458
0 3 14 0 0 8192 0 0 19 38 0 4
938 477
1100 477
1100 305
1123 305
0 2 15 0 0 4224 0 0 19 50 0 4
981 317
1077 317
1077 296
1123 296
0 1 16 0 0 8192 0 0 19 29 0 4
1004 159
1100 159
1100 287
1123 287
3 4 17 0 0 12416 0 20 27 0 0 4
492 398
532 398
532 319
852 319
2 3 18 0 0 4224 0 27 21 0 0 3
852 301
494 301
494 331
4 3 19 0 0 12416 0 28 22 0 0 6
852 177
762 177
762 237
496 237
496 270
493 270
2 3 20 0 0 4224 0 28 23 0 0 2
852 159
492 159
4 3 13 0 0 12416 0 26 13 0 0 4
847 476
618 476
618 492
307 492
3 1 21 0 0 12416 0 15 20 0 0 4
243 405
246 405
246 389
447 389
1 2 22 0 0 4224 0 21 11 0 0 2
449 322
357 322
3 1 23 0 0 12416 0 16 11 0 0 4
241 339
245 339
245 322
321 322
2 0 16 0 0 0 0 14 0 0 29 2
187 469
143 469
2 0 16 0 0 0 0 15 0 0 29 2
194 414
143 414
0 2 16 0 0 8320 0 0 16 53 0 5
1004 159
1004 617
143 617
143 348
192 348
3 1 24 0 0 8320 0 14 13 0 0 4
236 460
249 460
249 483
258 483
2 0 25 0 0 4096 0 13 0 0 36 2
258 501
169 501
3 1 26 0 0 4224 0 18 23 0 0 4
238 223
355 223
355 150
447 150
2 1 27 0 0 4224 0 12 22 0 0 2
359 261
448 261
3 1 28 0 0 12416 0 17 12 0 0 4
239 279
246 279
246 261
323 261
2 0 25 0 0 0 0 17 0 0 36 2
190 288
169 288
0 2 25 0 0 8320 0 0 18 52 0 5
957 299
957 596
169 596
169 232
189 232
2 0 14 0 0 0 0 22 0 0 38 2
448 279
380 279
0 2 14 0 0 8320 0 0 23 44 0 5
938 475
938 574
380 574
380 168
447 168
0 2 29 0 0 4096 0 0 20 40 0 2
401 407
447 407
0 2 29 0 0 8320 0 0 21 45 0 5
910 457
910 553
401 553
401 340
449 340
1 1 3 0 0 0 0 2 18 0 0 4
43 305
62 305
62 214
189 214
0 3 11 0 0 4096 0 0 26 48 0 3
807 305
807 467
841 467
4 1 30 0 0 8320 0 19 33 0 0 3
1168 296
1200 296
1200 160
1 6 14 0 0 0 0 24 26 0 0 4
936 431
938 431
938 476
901 476
7 1 29 0 0 0 0 26 25 0 0 3
895 458
910 458
910 429
5 0 31 0 0 8192 0 26 0 0 49 3
871 506
871 521
783 521
5 0 31 0 0 8192 0 27 0 0 49 3
876 349
876 355
783 355
0 3 11 0 0 4224 0 0 27 55 0 4
358 103
807 103
807 310
846 310
5 1 31 0 0 16512 0 28 3 0 0 5
876 207
876 210
783 210
783 523
41 523
6 1 15 0 0 0 0 27 29 0 0 3
906 319
981 319
981 262
6 1 32 0 0 4224 0 28 30 0 0 3
906 177
1027 177
1027 120
7 1 25 0 0 0 0 27 31 0 0 3
900 301
957 301
957 262
7 1 16 0 0 0 0 28 32 0 0 4
900 159
1006 159
1006 120
1005 120
0 1 10 0 0 0 0 0 28 0 0 4
875 123
875 126
876 126
876 132
6 1 11 0 0 0 0 38 34 0 0 3
251 103
359 103
359 70
0 1 2 0 0 4224 0 0 35 1 0 4
227 66
8 66
8 121
18 121
1 2 33 0 0 4224 0 4 38 0 0 4
59 88
188 88
188 103
203 103
4 1 34 0 0 4224 0 38 36 0 0 2
227 151
227 159
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
