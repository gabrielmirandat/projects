* C:\Users\Marina\Desktop\EXP6ABODE.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 27 12:56:51 2015



** Analysis setup **
.ac DEC 101 1K 100K


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EXP6ABODE.net"
.INC "EXP6ABODE.als"


.probe


.END
