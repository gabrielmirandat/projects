CircuitMaker Text
5.6
Probes: 3
ra[i]
Transient Analysis
0 420 165 65280
rd[i]
Transient Analysis
1 641 188 65535
rc[i]
Transient Analysis
2 638 274 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 120 30 100 10
321 166 1336 703
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 1 1 1
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
489 262 1504 530
1083744434 0
0
6 Title:
5 Name:
0
0
0
8
9 V Source~
197 363 232 0 2 5
0 5 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
5130 0 0
2
5.89725e-315 5.26354e-315
0
7 Ground~
168 446 324 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
5.89725e-315 0
0
9 Resistor~
219 437 164 0 2 5
0 5 6
0
0 0 880 0
4 2011
-14 -14 14 -6
2 Ra
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3124 0 0
2
5.89725e-315 5.37752e-315
0
9 Resistor~
219 553 203 0 2 5
0 4 6
0
0 0 880 90
4 1035
1 0 29 8
2 Rb
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
5.89725e-315 5.36716e-315
0
9 Resistor~
219 640 202 0 2 5
0 3 6
0
0 0 880 90
4 4700
3 0 31 8
2 Rd
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8157 0 0
2
5.89725e-315 5.3568e-315
0
9 Resistor~
219 601 248 0 2 5
0 3 4
0
0 0 880 180
3 100
-10 -14 11 -6
2 Rf
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5572 0 0
2
5.89725e-315 5.34643e-315
0
9 Resistor~
219 554 287 0 3 5
0 2 4 -1
0
0 0 880 90
4 4700
1 0 29 8
2 Re
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
5.89725e-315 5.32571e-315
0
9 Resistor~
219 640 289 0 3 5
0 2 3 -1
0
0 0 880 90
4 1035
1 0 29 8
2 Rc
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7361 0 0
2
5.89725e-315 5.30499e-315
0
10
1 0 2 0 0 4096 0 7 0 0 2 2
554 305
554 318
1 1 2 0 0 4224 0 2 8 0 0 3
446 318
640 318
640 307
2 1 2 0 0 0 0 1 2 0 0 3
363 253
363 318
446 318
1 0 3 0 0 4096 0 6 0 0 5 2
619 248
640 248
1 2 3 0 0 4224 0 5 8 0 0 2
640 220
640 271
2 0 4 0 0 4096 0 6 0 0 7 2
583 248
554 248
1 2 4 0 0 8320 0 4 7 0 0 3
553 221
554 221
554 269
2 0 6 0 0 4096 0 4 0 0 9 2
553 185
553 164
2 2 6 0 0 4224 0 3 5 0 0 3
455 164
640 164
640 184
1 1 5 0 0 8320 0 1 3 0 0 3
363 211
363 164
419 164
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
640 225 659 241
640 225 659 241
2 v4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
554 223 573 239
554 223 573 239
2 v3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
512 302 531 318
512 302 531 318
2 v0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
363 168 382 184
363 168 382 184
2 v1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
573 148 592 164
573 148 592 164
2 v2
0
17 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
