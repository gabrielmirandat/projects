CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 120 308 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
42179.7 0
0
13 Logic Switch~
5 121 240 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
317 0 0
2
42179.7 0
0
13 Logic Switch~
5 123 173 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3108 0 0
2
42179.7 0
0
13 Logic Switch~
5 125 105 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4299 0 0
2
42179.7 0
0
13 Logic Switch~
5 117 396 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 E1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
42179.7 0
0
13 Logic Switch~
5 118 478 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 E2
-4 -28 10 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7876 0 0
2
42179.7 0
0
14 Logic Display~
6 862 155 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
42179.7 0
0
5 4012~
219 726 208 0 5 22
0 6 5 4 3 2
0
0 0 624 0
4 4012
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 4 0
1 U
9172 0 0
2
42179.7 0
0
9 Inverter~
13 233 478 0 2 22
0 7 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7100 0 0
2
42179.7 0
0
9 Inverter~
13 233 396 0 2 22
0 8 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3820 0 0
2
42179.7 0
0
10 3-In NAND~
219 507 317 0 4 22
0 11 8 7 3
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
7678 0 0
2
42179.7 0
0
10 3-In NAND~
219 504 249 0 4 22
0 12 8 9 4
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 1 0
1 U
961 0 0
2
42179.7 0
0
10 3-In NAND~
219 505 182 0 4 22
0 13 10 7 5
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
3178 0 0
2
42179.7 0
0
10 3-In NAND~
219 506 114 0 4 22
0 14 10 9 6
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
3409 0 0
2
42179.7 0
0
19
5 1 2 0 0 4224 0 8 7 0 0 3
753 208
862 208
862 173
4 4 3 0 0 4224 0 11 8 0 0 4
534 317
682 317
682 222
702 222
4 3 4 0 0 4224 0 12 8 0 0 4
531 249
648 249
648 213
702 213
4 2 5 0 0 4224 0 13 8 0 0 4
532 182
649 182
649 204
702 204
4 1 6 0 0 4224 0 14 8 0 0 4
533 114
682 114
682 195
702 195
3 0 7 0 0 4096 0 11 0 0 10 2
483 326
448 326
2 0 8 0 0 4096 0 11 0 0 9 2
483 317
395 317
3 0 9 0 0 4096 0 12 0 0 12 2
480 258
289 258
0 2 8 0 0 8320 0 0 12 15 0 5
195 396
195 430
395 430
395 249
480 249
0 3 7 0 0 12416 0 0 13 14 0 5
195 478
195 516
448 516
448 191
481 191
2 0 10 0 0 4096 0 13 0 0 13 2
481 182
269 182
2 3 9 0 0 8320 0 9 14 0 0 4
254 478
289 478
289 123
482 123
2 2 10 0 0 8320 0 10 14 0 0 4
254 396
269 396
269 114
482 114
1 1 7 0 0 0 0 6 9 0 0 2
130 478
218 478
1 1 8 0 0 0 0 5 10 0 0 2
129 396
218 396
1 1 11 0 0 4224 0 1 11 0 0 2
132 308
483 308
1 1 12 0 0 4224 0 2 12 0 0 2
133 240
480 240
1 1 13 0 0 4224 0 3 13 0 0 2
135 173
481 173
1 1 14 0 0 4224 0 4 14 0 0 2
137 105
482 105
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
