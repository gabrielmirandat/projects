CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
43032754 0
0
6 Title:
5 Name:
0
0
0
61
13 Logic Switch~
5 44 502 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
5 NSCAR
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
42291 0
0
13 Logic Switch~
5 44 543 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 EWCAR
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
42291 1
0
7 Ground~
168 140 366 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
42291 2
0
7 Pulser~
4 324 168 0 10 12
0 82 83 12 84 0 0 5 5 5
7
0
0 0 4656 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3421 0 0
2
42291 3
0
10 StopLight~
181 1122 503 0 12 13
0 7 6 3 0 0 0 0 0 0
0 0 1
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM2
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
8157 0 0
2
42291 4
0
10 StopLight~
181 1120 401 0 10 13
0 8 5 4 0 0 0 0 0 0
1
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM1
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 1 0 0 0
3 SEM
5572 0 0
2
42291 5
0
9 Inverter~
13 950 571 0 2 22
0 15 4
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U16D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
8901 0 0
2
42291 6
0
9 Inverter~
13 951 528 0 2 22
0 13 3
0
0 0 624 0
5 74F04
-50 -22 -15 -14
4 U16C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
7361 0 0
2
42291 7
0
10 2-In NAND~
219 956 446 0 3 22
0 17 11 5
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4747 0 0
2
42291 8
0
10 2-In NAND~
219 957 489 0 3 22
0 14 16 6
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
972 0 0
2
42291 9
0
2 +V
167 919 266 0 1 3
0 20
0
0 0 54256 0
3 10V
29 -11 50 -3
2 V8
13 -11 27 -3
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
42291 10
0
10 8-In NAND~
219 957 392 0 9 19
0 20 20 20 19 18 17 11 15 7
0
0 0 624 0
6 74LS30
-21 -24 21 -16
3 U20
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
42291 11
0
10 8-In NAND~
219 957 315 0 9 19
0 20 20 20 19 16 14 13 18 8
0
0 0 624 0
6 74LS30
-21 -24 21 -16
3 U19
-12 -44 9 -36
0
15 DVCC=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 3 4 5 6 11 12 8
1 2 3 4 5 6 11 12 8 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
42291 12
0
7 Ground~
168 718 596 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
42291 13
0
2 +V
167 744 597 0 1 3
0 26
0
0 0 54256 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
42291 14
0
7 74LS138
19 790 535 0 14 29
0 23 22 21 26 2 2 19 16 14
13 18 17 11 15
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
3 U18
-11 -71 10 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
42291 15
0
7 Pulser~
4 67 411 0 10 12
0 85 86 27 87 0 0 5 5 5
7
0
0 0 4656 0
0
2 V2
-8 22 6 30
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5616 0 0
2
42291 16
0
2 +V
167 592 474 0 1 3
0 28
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
42291 17
0
7 Ground~
168 452 479 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
42291 18
0
9 Inverter~
13 602 505 0 2 22
0 25 24
0
0 0 624 180
5 74F04
13 -17 48 -9
4 U16B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
3108 0 0
2
42291 19
0
9 3-In AND~
219 640 559 0 4 22
0 23 22 21 25
0
0 0 624 0
6 74LS11
-23 21 19 29
4 U15C
-14 32 14 40
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 10 0
1 U
4299 0 0
2
42291 20
0
7 74LS161
96 542 532 0 14 29
0 29 29 27 88 89 90 91 28 24
92 93 23 22 21
0
0 0 4848 0
8 74LS161A
-27 -71 29 -63
3 U17
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
42291 21
0
8 2-In OR~
219 285 534 0 3 22
0 9 31 37
0
0 0 624 0
6 74LS32
5 -30 47 -22
4 U14B
-26 -29 2 -21
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
7876 0 0
2
42291 22
0
8 2-In OR~
219 285 570 0 3 22
0 9 30 36
0
0 0 624 0
6 74LS32
5 19 47 27
4 U14A
-23 20 5 28
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
6369 0 0
2
42291 23
0
2 +V
167 343 602 0 1 3
0 38
0
0 0 54256 180
3 10V
9 -3 30 5
2 V5
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9172 0 0
2
42291 24
0
7 74LS151
20 399 534 0 14 29
0 38 38 38 37 38 38 38 36 2
23 22 21 29 94
0
0 0 4848 0
7 74LS151
-24 -72 25 -64
3 U13
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7100 0 0
2
42291 25
0
9 Inverter~
13 260 287 0 2 22
0 77 9
0
0 0 624 270
5 74F04
-18 -19 17 -11
4 U16A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
3820 0 0
2
42291 26
0
9 3-In AND~
219 212 579 0 4 22
0 35 34 10 30
0
0 0 624 0
6 74LS11
-47 17 -5 25
4 U15B
2 17 30 25
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 10 0
1 U
7678 0 0
2
42291 27
0
9 3-In AND~
219 212 543 0 4 22
0 32 33 10 31
0
0 0 624 0
6 74LS11
-40 -26 2 -18
4 U15A
3 -26 31 -18
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 10 0
1 U
961 0 0
2
42291 28
0
9 Inverter~
13 95 522 0 2 22
0 34 32
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3178 0 0
2
42291 29
0
9 Inverter~
13 96 471 0 2 22
0 33 35
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3409 0 0
2
42291 30
0
2 +V
167 79 164 0 1 3
0 39
0
0 0 54256 180
3 10V
6 -2 27 6
2 V1
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
42291 31
0
9 4-In AND~
219 468 244 0 5 22
0 53 56 52 54 43
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U11A
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
8885 0 0
2
42291 32
0
9 Inverter~
13 388 218 0 2 22
0 55 53
0
0 0 624 0
5 74F04
-18 -30 17 -22
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3780 0 0
2
42291 33
0
9 Inverter~
13 389 252 0 2 22
0 57 52
0
0 0 624 0
5 74F04
13 -17 48 -9
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
9265 0 0
2
42291 34
0
9 Inverter~
13 387 340 0 2 22
0 51 46
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
9442 0 0
2
42291 35
0
9 Inverter~
13 388 302 0 2 22
0 49 47
0
0 0 624 0
5 74F04
-18 -30 17 -22
4 U10B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
9424 0 0
2
42291 36
0
9 4-In AND~
219 468 328 0 5 22
0 47 44 46 45 42
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 U11B
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
9968 0 0
2
42291 37
0
9 Inverter~
13 354 359 0 2 22
0 48 45
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
9281 0 0
2
42291 38
0
9 Inverter~
13 353 322 0 2 22
0 50 44
0
0 0 624 0
5 74F04
13 -17 48 -9
4 U10D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
8464 0 0
2
42291 39
0
9 2-In AND~
219 536 274 0 3 22
0 43 42 40
0
0 0 624 0
6 74LS08
-24 -36 18 -28
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
7168 0 0
2
42291 40
0
6 74LS48
188 1022 79 0 14 29
0 55 56 57 54 95 96 65 64 63
62 61 60 59 97
0
0 0 4848 0
6 74LS48
-21 -76 21 -68
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3171 0 0
2
42291 41
0
9 Inverter~
13 929 148 0 2 22
0 56 66
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U7C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
4139 0 0
2
42291 42
0
9 Inverter~
13 942 180 0 2 22
0 57 58
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U7B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
6435 0 0
2
42291 43
0
9 Inverter~
13 694 146 0 2 22
0 49 67
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U7F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
5283 0 0
2
42291 44
0
9 Inverter~
13 718 144 0 2 22
0 50 68
0
0 0 624 270
5 74F04
-18 -19 17 -11
3 U7E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
6874 0 0
2
42291 45
0
6 74LS48
188 814 78 0 14 29
0 49 50 51 48 98 99 75 74 73
72 71 70 69 100
0
0 0 4848 0
6 74LS48
-21 -76 21 -68
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5305 0 0
2
42291 46
0
10 4-In NAND~
219 617 94 0 5 22
0 54 58 66 55 76
0
0 0 624 180
6 74LS20
-21 -40 21 -32
3 U5A
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 1 0
1 U
34 0 0
2
42291 47
0
9 CC 7-Seg~
183 88 244 0 12 19
10 69 70 71 72 73 74 75 2 2
0 1 1
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP2
34 -4 69 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
969 0 0
2
42291 48
0
9 CC 7-Seg~
183 193 243 0 16 19
10 59 60 61 62 63 64 65 2 2
1 1 0 1 1 0 1
0
0 0 21088 0
7 AMBERCC
-77 -28 -28 -20
5 DISP1
-70 -15 -35 -7
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
8402 0 0
2
42291 49
0
7 74LS160
124 145 139 0 14 29
0 39 39 76 39 101 102 103 104 78
105 49 50 51 48
0
0 0 4848 0
8 74LS160A
-25 -61 31 -53
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3751 0 0
2
5.89727e-315 0
0
10 4-In NAND~
219 277 112 0 5 22
0 48 51 68 67 77
0
0 0 624 180
6 74LS20
-21 -40 21 -32
3 U5B
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
4292 0 0
2
5.89727e-315 5.26354e-315
0
14 Logic Display~
6 825 288 0 1 2
10 9
0
0 0 53856 0
6 100MEG
16 1 58 9
6 TMLONG
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.89727e-315 5.30499e-315
0
2 +V
167 612 200 0 1 3
0 41
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
34 0 0
2
5.89727e-315 5.32571e-315
0
14 Logic Display~
6 749 287 0 1 2
10 10
0
0 0 53856 0
6 100MEG
16 1 58 9
7 TMSHORT
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
5.89727e-315 5.34643e-315
0
10 2-In NAND~
219 264 38 0 3 22
0 8 7 80
0
0 0 624 0
4 7400
-15 -36 13 -28
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
319 0 0
2
5.89727e-315 5.3568e-315
0
9 2-In AND~
219 543 85 0 3 22
0 76 80 79
0
0 0 624 180
6 74LS08
-24 -36 18 -28
3 U9B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3976 0 0
2
5.89727e-315 5.36716e-315
0
9 2-In AND~
219 222 103 0 3 22
0 77 80 78
0
0 0 624 180
6 74LS08
-24 -36 18 -28
3 U9A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7634 0 0
2
5.89727e-315 5.37752e-315
0
7 74LS163
126 462 121 0 14 29
0 81 81 12 81 106 107 108 109 79
110 55 56 57 54
0
0 0 4848 0
8 74LS163A
-28 -62 28 -54
2 U2
-8 -52 6 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
523 0 0
2
5.89727e-315 5.38788e-315
0
5 7474~
219 612 292 0 6 22
0 41 41 40 78 111 10
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U8A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
6748 0 0
2
42291 50
0
2 +V
167 418 77 0 1 3
0 81
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6901 0 0
2
42291 51
0
192
2 0 11 0 0 4096 0 9 0 0 25 2
932 455
887 455
8 0 2 0 0 8192 0 49 0 0 5 3
109 280
109 299
129 299
8 0 2 0 0 8192 0 50 0 0 4 3
214 279
214 299
242 299
1 9 2 0 0 8320 0 3 50 0 0 4
140 360
242 360
242 201
193 201
9 1 2 0 0 0 0 49 3 0 0 4
88 202
129 202
129 360
140 360
3 3 12 0 0 8320 0 4 59 0 0 4
348 159
385 159
385 112
430 112
3 2 6 0 0 12416 0 10 5 0 0 4
984 489
1025 489
1025 503
1106 503
0 1 7 0 0 8320 0 0 5 13 0 4
991 392
1074 392
1074 489
1106 489
0 1 8 0 0 4224 0 0 6 14 0 4
994 315
1084 315
1084 387
1104 387
2 1 7 0 0 0 0 56 0 0 12 2
240 47
164 47
1 0 8 0 0 0 0 56 0 0 12 2
240 29
164 29
7 0 1 0 0 4128 0 0 0 0 0 2
164 20
164 55
9 1 7 0 0 0 0 12 0 0 15 4
984 392
991 392
991 349
1025 349
9 0 8 0 0 0 0 13 0 0 15 4
984 315
994 315
994 335
1025 335
7 0 1 0 0 4128 0 0 0 0 0 2
1025 322
1025 361
1 0 13 0 0 4096 0 8 0 0 36 2
936 528
863 528
1 0 14 0 0 4096 0 10 0 0 37 2
933 480
854 480
1 0 15 0 0 4096 0 7 0 0 24 2
935 571
894 571
2 0 16 0 0 4096 0 10 0 0 38 2
933 498
845 498
1 0 17 0 0 4096 0 9 0 0 26 2
932 437
879 437
2 3 4 0 0 16512 0 7 6 0 0 6
971 571
1062 571
1062 561
1087 561
1087 415
1104 415
2 3 3 0 0 4224 0 8 5 0 0 4
972 528
1062 528
1062 517
1106 517
3 2 5 0 0 4224 0 9 6 0 0 4
983 446
1059 446
1059 401
1104 401
14 8 15 0 0 8320 0 16 12 0 0 4
828 571
896 571
896 424
933 424
13 7 11 0 0 8320 0 16 12 0 0 4
828 562
887 562
887 415
933 415
12 6 17 0 0 8320 0 16 12 0 0 4
828 553
879 553
879 406
933 406
5 0 18 0 0 4096 0 12 0 0 35 2
933 397
871 397
4 0 19 0 0 4096 0 12 0 0 39 2
933 388
837 388
0 3 20 0 0 4096 0 0 12 30 0 2
919 379
933 379
0 2 20 0 0 0 0 0 12 31 0 5
919 370
919 379
919 379
919 370
933 370
0 1 20 0 0 4224 0 0 12 32 0 5
919 301
919 370
919 370
919 361
933 361
0 3 20 0 0 0 0 0 13 33 0 3
919 293
919 302
933 302
0 2 20 0 0 0 0 0 13 34 0 3
919 283
919 293
933 293
1 1 20 0 0 0 0 11 13 0 0 3
919 275
919 284
933 284
11 8 18 0 0 8320 0 16 13 0 0 4
828 544
871 544
871 347
933 347
10 7 13 0 0 8320 0 16 13 0 0 4
828 535
863 535
863 338
933 338
9 6 14 0 0 8320 0 16 13 0 0 4
828 526
854 526
854 329
933 329
8 5 16 0 0 8320 0 16 13 0 0 4
828 517
845 517
845 320
933 320
7 4 19 0 0 8320 0 16 13 0 0 4
828 508
837 508
837 311
933 311
0 12 21 0 0 8320 0 0 26 45 0 5
608 568
608 601
452 601
452 534
431 534
0 11 22 0 0 8320 0 0 26 44 0 5
601 559
601 593
461 593
461 525
431 525
0 10 23 0 0 8192 0 0 26 43 0 5
594 550
594 585
470 585
470 516
431 516
0 1 23 0 0 8320 0 0 16 57 0 5
594 550
594 522
719 522
719 508
758 508
0 2 22 0 0 0 0 0 16 58 0 5
601 559
601 530
727 530
727 517
758 517
0 3 21 0 0 0 0 0 16 56 0 5
608 568
608 539
735 539
735 526
758 526
2 9 24 0 0 12416 0 20 22 0 0 4
587 505
588 505
588 505
580 505
1 4 25 0 0 8320 0 20 21 0 0 4
623 505
673 505
673 559
661 559
0 5 2 0 0 0 0 0 16 49 0 3
718 572
718 562
752 562
1 6 2 0 0 0 0 14 16 0 0 3
718 590
718 571
752 571
1 4 26 0 0 4224 0 15 16 0 0 3
744 582
744 553
758 553
3 3 27 0 0 12416 0 22 17 0 0 4
510 514
494 514
494 402
91 402
8 1 28 0 0 8320 0 22 18 0 0 3
580 496
592 496
592 483
2 0 29 0 0 4096 0 22 0 0 54 2
510 505
475 505
13 1 29 0 0 8320 0 26 22 0 0 4
431 561
475 561
475 496
510 496
9 1 2 0 0 0 0 26 19 0 0 3
437 507
452 507
452 487
3 14 21 0 0 0 0 21 22 0 0 2
616 568
574 568
12 1 23 0 0 0 0 22 21 0 0 2
574 550
616 550
13 2 22 0 0 0 0 22 21 0 0 2
574 559
616 559
4 2 30 0 0 4224 0 28 24 0 0 2
233 579
272 579
4 2 31 0 0 4224 0 29 23 0 0 2
233 543
272 543
2 1 32 0 0 12416 0 30 29 0 0 4
116 522
138 522
138 534
188 534
0 2 33 0 0 4224 0 0 29 78 0 4
66 489
164 489
164 543
188 543
0 3 10 0 0 4096 0 0 28 64 0 3
173 552
173 588
188 588
0 3 10 0 0 8320 0 0 29 84 0 5
749 320
749 444
173 444
173 552
188 552
0 2 34 0 0 8320 0 0 28 77 0 3
66 543
66 579
188 579
2 1 35 0 0 8320 0 31 28 0 0 4
117 471
156 471
156 570
188 570
0 1 9 0 0 4096 0 0 24 68 0 3
263 523
263 561
272 561
0 1 9 0 0 4096 0 0 23 83 0 3
263 414
263 525
272 525
3 8 36 0 0 4224 0 24 26 0 0 2
318 570
367 570
3 4 37 0 0 4224 0 23 26 0 0 2
318 534
367 534
3 0 38 0 0 4096 0 26 0 0 73 2
367 525
343 525
2 0 38 0 0 0 0 26 0 0 73 2
367 516
343 516
0 1 38 0 0 4224 0 0 26 74 0 3
343 543
343 507
367 507
0 5 38 0 0 0 0 0 26 75 0 3
343 553
343 543
367 543
0 6 38 0 0 0 0 0 26 76 0 3
343 561
343 552
367 552
1 7 38 0 0 0 0 25 26 0 0 3
343 587
343 561
367 561
1 1 34 0 0 0 0 2 30 0 0 4
56 543
67 543
67 522
80 522
1 1 33 0 0 0 0 1 31 0 0 4
56 502
66 502
66 471
81 471
4 0 39 0 0 4096 0 51 0 0 81 2
107 139
79 139
2 0 39 0 0 4096 0 51 0 0 81 2
113 121
79 121
1 1 39 0 0 8320 0 51 32 0 0 3
113 112
79 112
79 149
3 3 40 0 0 4224 0 41 60 0 0 2
557 274
588 274
2 1 9 0 0 8320 0 27 53 0 0 4
263 305
263 415
825 415
825 306
6 1 10 0 0 0 0 60 55 0 0 5
636 256
675 256
675 320
749 320
749 305
2 0 41 0 0 12416 0 60 0 0 86 4
588 256
575 256
575 220
612 220
1 1 41 0 0 0 0 54 60 0 0 2
612 209
612 229
5 2 42 0 0 8320 0 38 41 0 0 4
489 328
502 328
502 283
512 283
5 1 43 0 0 8320 0 33 41 0 0 4
489 244
502 244
502 265
512 265
2 2 44 0 0 12416 0 40 38 0 0 4
374 322
381 322
381 324
444 324
2 4 45 0 0 4224 0 39 38 0 0 4
375 359
429 359
429 342
444 342
2 3 46 0 0 12416 0 36 38 0 0 4
408 340
425 340
425 333
444 333
2 1 47 0 0 12416 0 37 38 0 0 4
409 302
425 302
425 315
444 315
0 1 48 0 0 4096 0 0 39 97 0 4
301 346
333 346
333 359
339 359
3 1 49 0 0 12288 0 0 37 97 0 4
301 311
316 311
316 302
373 302
2 1 50 0 0 4096 0 0 40 97 0 2
301 322
338 322
1 1 51 0 0 12288 0 0 36 97 0 4
301 336
316 336
316 340
372 340
1 0 1 0 0 4128 0 0 0 0 0 2
301 302
301 351
2 3 52 0 0 12416 0 35 33 0 0 4
410 252
425 252
425 249
444 249
2 1 53 0 0 12416 0 34 33 0 0 4
409 218
425 218
425 231
444 231
0 4 54 0 0 12288 0 0 33 104 0 6
301 262
333 262
333 275
429 275
429 258
444 258
3 1 55 0 0 12288 0 0 34 104 0 4
301 227
316 227
316 218
373 218
2 2 56 0 0 4224 0 0 33 104 0 4
301 238
381 238
381 240
444 240
1 1 57 0 0 4096 0 0 35 104 0 2
301 252
374 252
4 0 1 0 0 32 0 0 0 0 0 2
301 218
301 267
2 1 58 0 0 4224 0 44 0 0 119 2
945 198
945 248
13 0 59 0 0 4096 0 42 0 0 113 2
1054 97
1093 97
12 1 60 0 0 4096 0 42 0 0 113 2
1054 88
1093 88
11 2 61 0 0 4096 0 42 0 0 113 2
1054 79
1093 79
10 3 62 0 0 4096 0 42 0 0 113 2
1054 70
1093 70
9 4 63 0 0 4096 0 42 0 0 113 2
1054 61
1093 61
8 5 64 0 0 4096 0 42 0 0 113 2
1054 52
1093 52
7 6 65 0 0 4096 0 42 0 0 113 2
1054 43
1093 43
6 0 1 0 0 4256 0 0 0 0 0 2
1093 35
1093 106
0 3 55 0 0 4224 0 0 0 120 119 4
920 43
920 239
925 239
925 248
2 2 66 0 0 4224 0 43 0 0 119 2
932 166
932 248
0 0 54 0 0 4224 0 0 0 123 119 4
975 70
975 207
958 207
958 248
0 1 57 0 0 4224 0 0 44 122 0 2
945 61
945 162
0 1 56 0 0 0 0 0 43 121 0 2
932 52
932 130
5 0 1 0 0 32 0 0 0 0 0 2
915 248
969 248
3 1 55 0 0 0 0 0 42 124 0 2
910 43
990 43
2 2 56 0 0 0 0 0 42 124 0 2
910 52
990 52
1 3 57 0 0 0 0 0 42 124 0 2
910 61
990 61
0 4 54 0 0 0 0 0 42 124 0 2
910 70
990 70
4 0 1 0 0 32 0 0 0 0 0 2
910 26
910 75
2 3 67 0 0 4224 0 45 0 0 139 4
697 164
697 219
719 219
719 247
2 2 68 0 0 4224 0 46 0 0 139 4
721 162
721 208
728 208
728 247
0 1 49 0 0 4096 0 0 45 140 0 4
715 42
715 105
697 105
697 128
1 0 50 0 0 4096 0 46 0 0 141 2
721 126
721 51
13 0 69 0 0 4096 0 47 0 0 136 2
846 96
885 96
12 1 70 0 0 4096 0 47 0 0 136 2
846 87
885 87
11 2 71 0 0 4096 0 47 0 0 136 2
846 78
885 78
10 3 72 0 0 4096 0 47 0 0 136 2
846 69
885 69
9 4 73 0 0 4096 0 47 0 0 136 2
846 60
885 60
8 5 74 0 0 4096 0 47 0 0 136 2
846 51
885 51
7 6 75 0 0 4096 0 47 0 0 136 2
846 42
885 42
3 0 1 0 0 32 0 0 0 0 0 2
885 34
885 105
0 0 48 0 0 4224 0 0 0 143 139 2
748 69
748 247
1 0 51 0 0 4224 0 0 0 139 142 2
735 247
735 60
2 0 1 0 0 32 0 0 0 0 0 2
705 247
759 247
3 1 49 0 0 4224 0 0 47 144 0 2
700 42
782 42
2 2 50 0 0 4224 0 0 47 144 0 2
700 51
782 51
1 3 51 0 0 0 0 0 47 144 0 2
700 60
782 60
0 4 48 0 0 0 0 0 47 144 0 2
700 69
782 69
1 0 1 0 0 32 0 0 0 0 0 2
700 25
700 74
5 0 76 0 0 4096 0 48 0 0 182 2
590 94
568 94
1 0 54 0 0 0 0 48 0 0 150 2
641 107
671 107
4 3 55 0 0 0 0 48 0 0 150 2
641 80
671 80
2 1 58 0 0 0 0 48 0 0 150 2
641 98
671 98
3 2 66 0 0 0 0 48 0 0 150 2
641 89
671 89
5 0 1 0 0 32 0 0 0 0 0 2
671 64
671 120
1 0 59 0 0 4224 0 50 0 0 158 2
172 279
172 325
2 1 60 0 0 4224 0 50 0 0 158 2
178 279
178 325
3 2 61 0 0 4224 0 50 0 0 158 2
184 279
184 325
4 3 62 0 0 4224 0 50 0 0 158 2
190 279
190 325
5 4 63 0 0 4224 0 50 0 0 158 2
196 279
196 325
6 5 64 0 0 4224 0 50 0 0 158 2
202 279
202 325
7 6 65 0 0 4224 0 50 0 0 158 2
208 279
208 325
6 0 1 0 0 32 0 0 0 0 0 2
163 325
227 325
1 0 69 0 0 4224 0 49 0 0 166 2
67 280
67 326
2 1 70 0 0 4224 0 49 0 0 166 2
73 280
73 326
3 2 71 0 0 4224 0 49 0 0 166 2
79 280
79 326
4 3 72 0 0 4224 0 49 0 0 166 2
85 280
85 326
5 4 73 0 0 4224 0 49 0 0 166 2
91 280
91 326
6 5 74 0 0 4224 0 49 0 0 166 2
97 280
97 326
7 6 75 0 0 4224 0 49 0 0 166 2
103 280
103 326
3 0 1 0 0 32 0 0 0 0 0 2
58 326
122 326
1 0 48 0 0 0 0 52 0 0 171 2
301 125
334 125
2 1 51 0 0 0 0 52 0 0 171 2
301 116
334 116
3 2 68 0 0 0 0 52 0 0 171 2
301 107
334 107
4 3 67 0 0 0 0 52 0 0 171 2
301 98
334 98
2 0 1 0 0 32 0 0 0 0 0 2
334 82
334 138
0 1 77 0 0 12416 0 0 27 178 0 4
245 112
245 150
263 150
263 269
0 4 78 0 0 16512 0 0 60 175 0 6
183 103
183 70
48 70
48 387
612 387
612 304
9 3 79 0 0 8320 0 59 57 0 0 4
500 94
508 94
508 85
516 85
9 3 78 0 0 0 0 51 58 0 0 3
183 112
183 103
195 103
0 2 80 0 0 4224 0 0 57 177 0 4
308 38
587 38
587 76
561 76
3 2 80 0 0 0 0 56 58 0 0 6
291 38
309 38
309 71
257 71
257 94
240 94
5 1 77 0 0 0 0 52 58 0 0 2
250 112
240 112
1 0 81 0 0 4096 0 59 0 0 181 2
430 94
418 94
2 0 81 0 0 0 0 59 0 0 181 2
430 103
418 103
1 4 81 0 0 4224 0 61 59 0 0 3
418 86
418 121
424 121
1 3 76 0 0 12416 0 57 51 0 0 6
561 94
569 94
569 196
94 196
94 130
113 130
11 3 55 0 0 0 0 59 0 0 187 2
494 130
538 130
12 2 56 0 0 0 0 59 0 0 187 2
494 139
538 139
13 1 57 0 0 0 0 59 0 0 187 2
494 148
538 148
14 0 54 0 0 0 0 59 0 0 187 2
494 157
538 157
4 0 1 0 0 32 0 0 0 0 0 2
538 116
538 165
11 3 49 0 0 0 0 51 0 0 192 2
177 148
220 148
12 2 50 0 0 0 0 51 0 0 192 2
177 157
220 157
13 1 51 0 0 0 0 51 0 0 192 2
177 166
220 166
14 0 48 0 0 0 0 51 0 0 192 2
177 175
220 175
1 0 1 0 0 32 0 0 0 0 0 2
220 134
220 183
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
988 512 1047 528
988 512 1047 528
7 EWGREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
989 555 1048 571
989 555 1048 571
7 NSGREEN
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 8
986 430 1053 446
986 430 1053 446
8 NSYELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 8
991 473 1058 489
991 473 1058 489
8 EWYELLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
1001 376 1044 392
1001 376 1044 392
5 EWRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
992 299 1035 315
992 299 1035 315
5 NSRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
185 31 228 47
185 31 228 47
5 EWRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
188 13 231 29
188 13 231 29
5 NSRED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 6
679 399 730 415
679 399 730 415
6 TMLONG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 7
676 304 735 320
676 304 735 320
7 TMSHORT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
