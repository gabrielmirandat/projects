* C:\Users\Marina\Desktop\EXP6A.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 27 13:09:29 2015



** Analysis setup **
.tran 1ns 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EXP6A.net"
.INC "EXP6A.als"


.probe


.END
