* C:\Users\gabriel\Dropbox\SEMESTRE6\7.CE2Lab\projects\proj6\simu\EXP6.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 18 19:16:31 2016



** Analysis setup **
.tran 1ns 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EXP6.net"
.INC "EXP6.als"


.probe


.END
