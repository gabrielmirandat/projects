CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Program Files\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
43024402 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 433 161 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 G
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89713e-315 0
0
13 Logic Switch~
5 434 118 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 F
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89713e-315 5.26354e-315
0
13 Logic Switch~
5 435 75 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 E
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89713e-315 5.30499e-315
0
13 Logic Switch~
5 40 226 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89713e-315 5.32571e-315
0
13 Logic Switch~
5 36 371 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
42179.7 0
0
13 Logic Switch~
5 37 324 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
42179.7 1
0
13 Logic Switch~
5 39 275 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
42179.7 2
0
14 Logic Display~
6 722 234 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
42179.7 3
0
10 2-In NAND~
219 348 236 0 3 22
0 8 7 6
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
4747 0 0
2
42179.7 4
0
10 2-In NAND~
219 346 283 0 3 22
0 5 5 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
972 0 0
2
42179.7 5
0
10 2-In NAND~
219 345 190 0 3 22
0 11 10 9
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3472 0 0
2
42179.7 6
0
2 +V
167 475 20 0 1 3
0 14
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
42179.7 7
0
7 Ground~
168 446 418 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
42179.7 8
0
7 Ground~
168 172 412 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
42179.7 9
0
10 2-In NAND~
219 345 328 0 3 22
0 8 12 13
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3835 0 0
2
42179.7 10
0
7 74LS154
95 247 265 0 22 45
0 2 2 18 21 20 19 8 22 23
24 11 10 7 25 5 26 27 28 29
30 31 12
0
0 0 4848 0
6 74F154
-21 -87 21 -79
2 U2
-7 -88 7 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
42179.7 11
0
7 74LS151
20 534 262 0 14 29
0 2 9 2 6 14 4 13 2 2
17 16 15 3 32
0
0 0 4848 0
6 74F151
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
42179.7 12
0
27
9 0 2 0 0 8192 0 17 0 0 18 4
572 235
572 192
446 192
446 235
13 1 3 0 0 4224 0 17 8 0 0 3
566 289
722 289
722 252
3 6 4 0 0 12416 0 10 17 0 0 4
373 283
419 283
419 280
502 280
0 2 5 0 0 8192 0 0 10 5 0 3
299 274
299 292
322 292
15 1 5 0 0 4224 0 16 10 0 0 2
285 274
322 274
3 4 6 0 0 12416 0 9 17 0 0 4
375 236
393 236
393 262
502 262
13 2 7 0 0 4224 0 16 9 0 0 4
285 256
316 256
316 245
324 245
0 1 8 0 0 4096 0 0 9 13 0 2
310 227
324 227
2 3 9 0 0 4224 0 17 11 0 0 4
502 244
404 244
404 190
372 190
12 2 10 0 0 8320 0 16 11 0 0 6
285 247
304 247
304 191
317 191
317 199
321 199
11 1 11 0 0 8320 0 16 11 0 0 4
285 238
298 238
298 181
321 181
22 2 12 0 0 4224 0 16 15 0 0 2
285 337
321 337
7 1 8 0 0 8320 0 16 15 0 0 4
285 202
310 202
310 319
321 319
7 3 13 0 0 8320 0 17 15 0 0 3
502 289
502 328
372 328
5 1 14 0 0 8320 0 17 12 0 0 3
502 271
475 271
475 29
8 0 2 0 0 0 0 17 0 0 18 2
502 298
446 298
3 0 2 0 0 0 0 17 0 0 18 2
502 253
446 253
1 1 2 0 0 8320 0 17 13 0 0 3
502 235
446 235
446 412
2 0 2 0 0 0 0 16 0 0 20 2
209 256
172 256
1 1 2 0 0 0 0 16 14 0 0 3
209 247
172 247
172 406
1 12 15 0 0 4224 0 1 17 0 0 4
445 161
640 161
640 262
566 262
1 11 16 0 0 4224 0 2 17 0 0 4
446 118
616 118
616 253
566 253
1 10 17 0 0 8320 0 3 17 0 0 4
447 75
593 75
593 244
566 244
3 1 18 0 0 12416 0 16 4 0 0 4
215 283
142 283
142 226
52 226
6 1 19 0 0 12416 0 16 5 0 0 4
215 310
142 310
142 371
48 371
5 1 20 0 0 4224 0 16 6 0 0 4
215 301
94 301
94 324
49 324
4 1 21 0 0 4224 0 16 7 0 0 4
215 292
94 292
94 275
51 275
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
